library verilog;
use verilog.vl_types.all;
entity axi_interconnect_v1_06_a is
    generic(
        C_FAMILY        : string  := "rtl";
        C_NUM_SLAVE_PORTS: integer := 2;
        C_THREAD_ID_WIDTH: integer := 0;
        C_THREAD_ID_PORT_WIDTH: integer := 1;
        C_AXI_ADDR_WIDTH: integer := 32;
        C_S00_AXI_DATA_WIDTH: integer := 32;
        C_S01_AXI_DATA_WIDTH: integer := 32;
        C_S02_AXI_DATA_WIDTH: integer := 32;
        C_S03_AXI_DATA_WIDTH: integer := 32;
        C_S04_AXI_DATA_WIDTH: integer := 32;
        C_S05_AXI_DATA_WIDTH: integer := 32;
        C_S06_AXI_DATA_WIDTH: integer := 32;
        C_S07_AXI_DATA_WIDTH: integer := 32;
        C_S08_AXI_DATA_WIDTH: integer := 32;
        C_S09_AXI_DATA_WIDTH: integer := 32;
        C_S10_AXI_DATA_WIDTH: integer := 32;
        C_S11_AXI_DATA_WIDTH: integer := 32;
        C_S12_AXI_DATA_WIDTH: integer := 32;
        C_S13_AXI_DATA_WIDTH: integer := 32;
        C_S14_AXI_DATA_WIDTH: integer := 32;
        C_S15_AXI_DATA_WIDTH: integer := 32;
        C_M00_AXI_DATA_WIDTH: integer := 32;
        C_INTERCONNECT_DATA_WIDTH: integer := 32;
        C_S00_AXI_ACLK_RATIO: string  := "1:1";
        C_S01_AXI_ACLK_RATIO: string  := "1:1";
        C_S02_AXI_ACLK_RATIO: string  := "1:1";
        C_S03_AXI_ACLK_RATIO: string  := "1:1";
        C_S04_AXI_ACLK_RATIO: string  := "1:1";
        C_S05_AXI_ACLK_RATIO: string  := "1:1";
        C_S06_AXI_ACLK_RATIO: string  := "1:1";
        C_S07_AXI_ACLK_RATIO: string  := "1:1";
        C_S08_AXI_ACLK_RATIO: string  := "1:1";
        C_S09_AXI_ACLK_RATIO: string  := "1:1";
        C_S10_AXI_ACLK_RATIO: string  := "1:1";
        C_S11_AXI_ACLK_RATIO: string  := "1:1";
        C_S12_AXI_ACLK_RATIO: string  := "1:1";
        C_S13_AXI_ACLK_RATIO: string  := "1:1";
        C_S14_AXI_ACLK_RATIO: string  := "1:1";
        C_S15_AXI_ACLK_RATIO: string  := "1:1";
        C_S00_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S01_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S02_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S03_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S04_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S05_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S06_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S07_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S08_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S09_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S10_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S11_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S12_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S13_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S14_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S15_AXI_IS_ACLK_ASYNC: integer := 0;
        C_M00_AXI_ACLK_RATIO: string  := "1:1";
        C_M00_AXI_IS_ACLK_ASYNC: integer := 0;
        C_S00_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S01_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S02_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S03_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S04_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S05_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S06_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S07_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S08_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S09_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S10_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S11_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S12_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S13_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S14_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S15_AXI_READ_WRITE_SUPPORT: string  := "READ/WRITE";
        C_S00_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S01_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S02_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S03_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S04_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S05_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S06_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S07_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S08_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S09_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S10_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S11_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S12_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S13_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S14_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S15_AXI_WRITE_ACCEPTANCE: integer := 1;
        C_S00_AXI_READ_ACCEPTANCE: integer := 1;
        C_S01_AXI_READ_ACCEPTANCE: integer := 1;
        C_S02_AXI_READ_ACCEPTANCE: integer := 1;
        C_S03_AXI_READ_ACCEPTANCE: integer := 1;
        C_S04_AXI_READ_ACCEPTANCE: integer := 1;
        C_S05_AXI_READ_ACCEPTANCE: integer := 1;
        C_S06_AXI_READ_ACCEPTANCE: integer := 1;
        C_S07_AXI_READ_ACCEPTANCE: integer := 1;
        C_S08_AXI_READ_ACCEPTANCE: integer := 1;
        C_S09_AXI_READ_ACCEPTANCE: integer := 1;
        C_S10_AXI_READ_ACCEPTANCE: integer := 1;
        C_S11_AXI_READ_ACCEPTANCE: integer := 1;
        C_S12_AXI_READ_ACCEPTANCE: integer := 1;
        C_S13_AXI_READ_ACCEPTANCE: integer := 1;
        C_S14_AXI_READ_ACCEPTANCE: integer := 1;
        C_S15_AXI_READ_ACCEPTANCE: integer := 1;
        C_M00_AXI_WRITE_ISSUING: integer := 1;
        C_M00_AXI_READ_ISSUING: integer := 1;
        C_S00_AXI_ARB_PRIORITY: integer := 0;
        C_S01_AXI_ARB_PRIORITY: integer := 0;
        C_S02_AXI_ARB_PRIORITY: integer := 0;
        C_S03_AXI_ARB_PRIORITY: integer := 0;
        C_S04_AXI_ARB_PRIORITY: integer := 0;
        C_S05_AXI_ARB_PRIORITY: integer := 0;
        C_S06_AXI_ARB_PRIORITY: integer := 0;
        C_S07_AXI_ARB_PRIORITY: integer := 0;
        C_S08_AXI_ARB_PRIORITY: integer := 0;
        C_S09_AXI_ARB_PRIORITY: integer := 0;
        C_S10_AXI_ARB_PRIORITY: integer := 0;
        C_S11_AXI_ARB_PRIORITY: integer := 0;
        C_S12_AXI_ARB_PRIORITY: integer := 0;
        C_S13_AXI_ARB_PRIORITY: integer := 0;
        C_S14_AXI_ARB_PRIORITY: integer := 0;
        C_S15_AXI_ARB_PRIORITY: integer := 0;
        C_S00_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S01_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S02_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S03_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S04_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S05_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S06_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S07_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S08_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S09_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S10_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S11_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S12_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S13_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S14_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S15_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_S00_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S01_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S02_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S03_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S04_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S05_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S06_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S07_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S08_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S09_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S10_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S11_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S12_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S13_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S14_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S15_AXI_READ_FIFO_DEPTH: integer := 0;
        C_M00_AXI_WRITE_FIFO_DEPTH: integer := 0;
        C_M00_AXI_READ_FIFO_DEPTH: integer := 0;
        C_S00_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S01_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S02_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S03_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S04_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S05_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S06_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S07_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S08_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S09_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S10_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S11_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S12_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S13_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S14_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S15_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_S00_AXI_READ_FIFO_DELAY: integer := 0;
        C_S01_AXI_READ_FIFO_DELAY: integer := 0;
        C_S02_AXI_READ_FIFO_DELAY: integer := 0;
        C_S03_AXI_READ_FIFO_DELAY: integer := 0;
        C_S04_AXI_READ_FIFO_DELAY: integer := 0;
        C_S05_AXI_READ_FIFO_DELAY: integer := 0;
        C_S06_AXI_READ_FIFO_DELAY: integer := 0;
        C_S07_AXI_READ_FIFO_DELAY: integer := 0;
        C_S08_AXI_READ_FIFO_DELAY: integer := 0;
        C_S09_AXI_READ_FIFO_DELAY: integer := 0;
        C_S10_AXI_READ_FIFO_DELAY: integer := 0;
        C_S11_AXI_READ_FIFO_DELAY: integer := 0;
        C_S12_AXI_READ_FIFO_DELAY: integer := 0;
        C_S13_AXI_READ_FIFO_DELAY: integer := 0;
        C_S14_AXI_READ_FIFO_DELAY: integer := 0;
        C_S15_AXI_READ_FIFO_DELAY: integer := 0;
        C_M00_AXI_WRITE_FIFO_DELAY: integer := 0;
        C_M00_AXI_READ_FIFO_DELAY: integer := 0;
        C_S00_AXI_REGISTER: integer := 0;
        C_S01_AXI_REGISTER: integer := 0;
        C_S02_AXI_REGISTER: integer := 0;
        C_S03_AXI_REGISTER: integer := 0;
        C_S04_AXI_REGISTER: integer := 0;
        C_S05_AXI_REGISTER: integer := 0;
        C_S06_AXI_REGISTER: integer := 0;
        C_S07_AXI_REGISTER: integer := 0;
        C_S08_AXI_REGISTER: integer := 0;
        C_S09_AXI_REGISTER: integer := 0;
        C_S10_AXI_REGISTER: integer := 0;
        C_S11_AXI_REGISTER: integer := 0;
        C_S12_AXI_REGISTER: integer := 0;
        C_S13_AXI_REGISTER: integer := 0;
        C_S14_AXI_REGISTER: integer := 0;
        C_S15_AXI_REGISTER: integer := 0;
        C_M00_AXI_REGISTER: integer := 0
    );
    port(
        INTERCONNECT_ACLK: in     vl_logic;
        INTERCONNECT_ARESETN: in     vl_logic;
        S00_AXI_ARESET_OUT_N: out    vl_logic;
        S00_AXI_ACLK    : in     vl_logic;
        S00_AXI_AWID    : in     vl_logic_vector;
        S00_AXI_AWADDR  : in     vl_logic_vector;
        S00_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S00_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S00_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S00_AXI_AWLOCK  : in     vl_logic;
        S00_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S00_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S00_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S00_AXI_AWVALID : in     vl_logic;
        S00_AXI_AWREADY : out    vl_logic;
        S00_AXI_WDATA   : in     vl_logic_vector;
        S00_AXI_WSTRB   : in     vl_logic_vector;
        S00_AXI_WLAST   : in     vl_logic;
        S00_AXI_WVALID  : in     vl_logic;
        S00_AXI_WREADY  : out    vl_logic;
        S00_AXI_BID     : out    vl_logic_vector;
        S00_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S00_AXI_BVALID  : out    vl_logic;
        S00_AXI_BREADY  : in     vl_logic;
        S00_AXI_ARID    : in     vl_logic_vector;
        S00_AXI_ARADDR  : in     vl_logic_vector;
        S00_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S00_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S00_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S00_AXI_ARLOCK  : in     vl_logic;
        S00_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S00_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S00_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S00_AXI_ARVALID : in     vl_logic;
        S00_AXI_ARREADY : out    vl_logic;
        S00_AXI_RID     : out    vl_logic_vector;
        S00_AXI_RDATA   : out    vl_logic_vector;
        S00_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S00_AXI_RLAST   : out    vl_logic;
        S00_AXI_RVALID  : out    vl_logic;
        S00_AXI_RREADY  : in     vl_logic;
        S01_AXI_ARESET_OUT_N: out    vl_logic;
        S01_AXI_ACLK    : in     vl_logic;
        S01_AXI_AWID    : in     vl_logic_vector;
        S01_AXI_AWADDR  : in     vl_logic_vector;
        S01_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S01_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S01_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S01_AXI_AWLOCK  : in     vl_logic;
        S01_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S01_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S01_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S01_AXI_AWVALID : in     vl_logic;
        S01_AXI_AWREADY : out    vl_logic;
        S01_AXI_WDATA   : in     vl_logic_vector;
        S01_AXI_WSTRB   : in     vl_logic_vector;
        S01_AXI_WLAST   : in     vl_logic;
        S01_AXI_WVALID  : in     vl_logic;
        S01_AXI_WREADY  : out    vl_logic;
        S01_AXI_BID     : out    vl_logic_vector;
        S01_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S01_AXI_BVALID  : out    vl_logic;
        S01_AXI_BREADY  : in     vl_logic;
        S01_AXI_ARID    : in     vl_logic_vector;
        S01_AXI_ARADDR  : in     vl_logic_vector;
        S01_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S01_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S01_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S01_AXI_ARLOCK  : in     vl_logic;
        S01_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S01_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S01_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S01_AXI_ARVALID : in     vl_logic;
        S01_AXI_ARREADY : out    vl_logic;
        S01_AXI_RID     : out    vl_logic_vector;
        S01_AXI_RDATA   : out    vl_logic_vector;
        S01_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S01_AXI_RLAST   : out    vl_logic;
        S01_AXI_RVALID  : out    vl_logic;
        S01_AXI_RREADY  : in     vl_logic;
        S02_AXI_ARESET_OUT_N: out    vl_logic;
        S02_AXI_ACLK    : in     vl_logic;
        S02_AXI_AWID    : in     vl_logic_vector;
        S02_AXI_AWADDR  : in     vl_logic_vector;
        S02_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S02_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S02_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S02_AXI_AWLOCK  : in     vl_logic;
        S02_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S02_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S02_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S02_AXI_AWVALID : in     vl_logic;
        S02_AXI_AWREADY : out    vl_logic;
        S02_AXI_WDATA   : in     vl_logic_vector;
        S02_AXI_WSTRB   : in     vl_logic_vector;
        S02_AXI_WLAST   : in     vl_logic;
        S02_AXI_WVALID  : in     vl_logic;
        S02_AXI_WREADY  : out    vl_logic;
        S02_AXI_BID     : out    vl_logic_vector;
        S02_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S02_AXI_BVALID  : out    vl_logic;
        S02_AXI_BREADY  : in     vl_logic;
        S02_AXI_ARID    : in     vl_logic_vector;
        S02_AXI_ARADDR  : in     vl_logic_vector;
        S02_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S02_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S02_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S02_AXI_ARLOCK  : in     vl_logic;
        S02_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S02_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S02_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S02_AXI_ARVALID : in     vl_logic;
        S02_AXI_ARREADY : out    vl_logic;
        S02_AXI_RID     : out    vl_logic_vector;
        S02_AXI_RDATA   : out    vl_logic_vector;
        S02_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S02_AXI_RLAST   : out    vl_logic;
        S02_AXI_RVALID  : out    vl_logic;
        S02_AXI_RREADY  : in     vl_logic;
        S03_AXI_ARESET_OUT_N: out    vl_logic;
        S03_AXI_ACLK    : in     vl_logic;
        S03_AXI_AWID    : in     vl_logic_vector;
        S03_AXI_AWADDR  : in     vl_logic_vector;
        S03_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S03_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S03_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S03_AXI_AWLOCK  : in     vl_logic;
        S03_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S03_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S03_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S03_AXI_AWVALID : in     vl_logic;
        S03_AXI_AWREADY : out    vl_logic;
        S03_AXI_WDATA   : in     vl_logic_vector;
        S03_AXI_WSTRB   : in     vl_logic_vector;
        S03_AXI_WLAST   : in     vl_logic;
        S03_AXI_WVALID  : in     vl_logic;
        S03_AXI_WREADY  : out    vl_logic;
        S03_AXI_BID     : out    vl_logic_vector;
        S03_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S03_AXI_BVALID  : out    vl_logic;
        S03_AXI_BREADY  : in     vl_logic;
        S03_AXI_ARID    : in     vl_logic_vector;
        S03_AXI_ARADDR  : in     vl_logic_vector;
        S03_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S03_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S03_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S03_AXI_ARLOCK  : in     vl_logic;
        S03_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S03_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S03_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S03_AXI_ARVALID : in     vl_logic;
        S03_AXI_ARREADY : out    vl_logic;
        S03_AXI_RID     : out    vl_logic_vector;
        S03_AXI_RDATA   : out    vl_logic_vector;
        S03_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S03_AXI_RLAST   : out    vl_logic;
        S03_AXI_RVALID  : out    vl_logic;
        S03_AXI_RREADY  : in     vl_logic;
        S04_AXI_ARESET_OUT_N: out    vl_logic;
        S04_AXI_ACLK    : in     vl_logic;
        S04_AXI_AWID    : in     vl_logic_vector;
        S04_AXI_AWADDR  : in     vl_logic_vector;
        S04_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S04_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S04_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S04_AXI_AWLOCK  : in     vl_logic;
        S04_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S04_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S04_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S04_AXI_AWVALID : in     vl_logic;
        S04_AXI_AWREADY : out    vl_logic;
        S04_AXI_WDATA   : in     vl_logic_vector;
        S04_AXI_WSTRB   : in     vl_logic_vector;
        S04_AXI_WLAST   : in     vl_logic;
        S04_AXI_WVALID  : in     vl_logic;
        S04_AXI_WREADY  : out    vl_logic;
        S04_AXI_BID     : out    vl_logic_vector;
        S04_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S04_AXI_BVALID  : out    vl_logic;
        S04_AXI_BREADY  : in     vl_logic;
        S04_AXI_ARID    : in     vl_logic_vector;
        S04_AXI_ARADDR  : in     vl_logic_vector;
        S04_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S04_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S04_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S04_AXI_ARLOCK  : in     vl_logic;
        S04_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S04_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S04_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S04_AXI_ARVALID : in     vl_logic;
        S04_AXI_ARREADY : out    vl_logic;
        S04_AXI_RID     : out    vl_logic_vector;
        S04_AXI_RDATA   : out    vl_logic_vector;
        S04_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S04_AXI_RLAST   : out    vl_logic;
        S04_AXI_RVALID  : out    vl_logic;
        S04_AXI_RREADY  : in     vl_logic;
        S05_AXI_ARESET_OUT_N: out    vl_logic;
        S05_AXI_ACLK    : in     vl_logic;
        S05_AXI_AWID    : in     vl_logic_vector;
        S05_AXI_AWADDR  : in     vl_logic_vector;
        S05_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S05_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S05_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S05_AXI_AWLOCK  : in     vl_logic;
        S05_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S05_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S05_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S05_AXI_AWVALID : in     vl_logic;
        S05_AXI_AWREADY : out    vl_logic;
        S05_AXI_WDATA   : in     vl_logic_vector;
        S05_AXI_WSTRB   : in     vl_logic_vector;
        S05_AXI_WLAST   : in     vl_logic;
        S05_AXI_WVALID  : in     vl_logic;
        S05_AXI_WREADY  : out    vl_logic;
        S05_AXI_BID     : out    vl_logic_vector;
        S05_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S05_AXI_BVALID  : out    vl_logic;
        S05_AXI_BREADY  : in     vl_logic;
        S05_AXI_ARID    : in     vl_logic_vector;
        S05_AXI_ARADDR  : in     vl_logic_vector;
        S05_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S05_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S05_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S05_AXI_ARLOCK  : in     vl_logic;
        S05_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S05_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S05_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S05_AXI_ARVALID : in     vl_logic;
        S05_AXI_ARREADY : out    vl_logic;
        S05_AXI_RID     : out    vl_logic_vector;
        S05_AXI_RDATA   : out    vl_logic_vector;
        S05_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S05_AXI_RLAST   : out    vl_logic;
        S05_AXI_RVALID  : out    vl_logic;
        S05_AXI_RREADY  : in     vl_logic;
        S06_AXI_ARESET_OUT_N: out    vl_logic;
        S06_AXI_ACLK    : in     vl_logic;
        S06_AXI_AWID    : in     vl_logic_vector;
        S06_AXI_AWADDR  : in     vl_logic_vector;
        S06_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S06_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S06_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S06_AXI_AWLOCK  : in     vl_logic;
        S06_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S06_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S06_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S06_AXI_AWVALID : in     vl_logic;
        S06_AXI_AWREADY : out    vl_logic;
        S06_AXI_WDATA   : in     vl_logic_vector;
        S06_AXI_WSTRB   : in     vl_logic_vector;
        S06_AXI_WLAST   : in     vl_logic;
        S06_AXI_WVALID  : in     vl_logic;
        S06_AXI_WREADY  : out    vl_logic;
        S06_AXI_BID     : out    vl_logic_vector;
        S06_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S06_AXI_BVALID  : out    vl_logic;
        S06_AXI_BREADY  : in     vl_logic;
        S06_AXI_ARID    : in     vl_logic_vector;
        S06_AXI_ARADDR  : in     vl_logic_vector;
        S06_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S06_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S06_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S06_AXI_ARLOCK  : in     vl_logic;
        S06_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S06_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S06_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S06_AXI_ARVALID : in     vl_logic;
        S06_AXI_ARREADY : out    vl_logic;
        S06_AXI_RID     : out    vl_logic_vector;
        S06_AXI_RDATA   : out    vl_logic_vector;
        S06_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S06_AXI_RLAST   : out    vl_logic;
        S06_AXI_RVALID  : out    vl_logic;
        S06_AXI_RREADY  : in     vl_logic;
        S07_AXI_ARESET_OUT_N: out    vl_logic;
        S07_AXI_ACLK    : in     vl_logic;
        S07_AXI_AWID    : in     vl_logic_vector;
        S07_AXI_AWADDR  : in     vl_logic_vector;
        S07_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S07_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S07_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S07_AXI_AWLOCK  : in     vl_logic;
        S07_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S07_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S07_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S07_AXI_AWVALID : in     vl_logic;
        S07_AXI_AWREADY : out    vl_logic;
        S07_AXI_WDATA   : in     vl_logic_vector;
        S07_AXI_WSTRB   : in     vl_logic_vector;
        S07_AXI_WLAST   : in     vl_logic;
        S07_AXI_WVALID  : in     vl_logic;
        S07_AXI_WREADY  : out    vl_logic;
        S07_AXI_BID     : out    vl_logic_vector;
        S07_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S07_AXI_BVALID  : out    vl_logic;
        S07_AXI_BREADY  : in     vl_logic;
        S07_AXI_ARID    : in     vl_logic_vector;
        S07_AXI_ARADDR  : in     vl_logic_vector;
        S07_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S07_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S07_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S07_AXI_ARLOCK  : in     vl_logic;
        S07_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S07_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S07_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S07_AXI_ARVALID : in     vl_logic;
        S07_AXI_ARREADY : out    vl_logic;
        S07_AXI_RID     : out    vl_logic_vector;
        S07_AXI_RDATA   : out    vl_logic_vector;
        S07_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S07_AXI_RLAST   : out    vl_logic;
        S07_AXI_RVALID  : out    vl_logic;
        S07_AXI_RREADY  : in     vl_logic;
        S08_AXI_ARESET_OUT_N: out    vl_logic;
        S08_AXI_ACLK    : in     vl_logic;
        S08_AXI_AWID    : in     vl_logic_vector;
        S08_AXI_AWADDR  : in     vl_logic_vector;
        S08_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S08_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S08_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S08_AXI_AWLOCK  : in     vl_logic;
        S08_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S08_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S08_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S08_AXI_AWVALID : in     vl_logic;
        S08_AXI_AWREADY : out    vl_logic;
        S08_AXI_WDATA   : in     vl_logic_vector;
        S08_AXI_WSTRB   : in     vl_logic_vector;
        S08_AXI_WLAST   : in     vl_logic;
        S08_AXI_WVALID  : in     vl_logic;
        S08_AXI_WREADY  : out    vl_logic;
        S08_AXI_BID     : out    vl_logic_vector;
        S08_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S08_AXI_BVALID  : out    vl_logic;
        S08_AXI_BREADY  : in     vl_logic;
        S08_AXI_ARID    : in     vl_logic_vector;
        S08_AXI_ARADDR  : in     vl_logic_vector;
        S08_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S08_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S08_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S08_AXI_ARLOCK  : in     vl_logic;
        S08_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S08_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S08_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S08_AXI_ARVALID : in     vl_logic;
        S08_AXI_ARREADY : out    vl_logic;
        S08_AXI_RID     : out    vl_logic_vector;
        S08_AXI_RDATA   : out    vl_logic_vector;
        S08_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S08_AXI_RLAST   : out    vl_logic;
        S08_AXI_RVALID  : out    vl_logic;
        S08_AXI_RREADY  : in     vl_logic;
        S09_AXI_ARESET_OUT_N: out    vl_logic;
        S09_AXI_ACLK    : in     vl_logic;
        S09_AXI_AWID    : in     vl_logic_vector;
        S09_AXI_AWADDR  : in     vl_logic_vector;
        S09_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S09_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S09_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S09_AXI_AWLOCK  : in     vl_logic;
        S09_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S09_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S09_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S09_AXI_AWVALID : in     vl_logic;
        S09_AXI_AWREADY : out    vl_logic;
        S09_AXI_WDATA   : in     vl_logic_vector;
        S09_AXI_WSTRB   : in     vl_logic_vector;
        S09_AXI_WLAST   : in     vl_logic;
        S09_AXI_WVALID  : in     vl_logic;
        S09_AXI_WREADY  : out    vl_logic;
        S09_AXI_BID     : out    vl_logic_vector;
        S09_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S09_AXI_BVALID  : out    vl_logic;
        S09_AXI_BREADY  : in     vl_logic;
        S09_AXI_ARID    : in     vl_logic_vector;
        S09_AXI_ARADDR  : in     vl_logic_vector;
        S09_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S09_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S09_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S09_AXI_ARLOCK  : in     vl_logic;
        S09_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S09_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S09_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S09_AXI_ARVALID : in     vl_logic;
        S09_AXI_ARREADY : out    vl_logic;
        S09_AXI_RID     : out    vl_logic_vector;
        S09_AXI_RDATA   : out    vl_logic_vector;
        S09_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S09_AXI_RLAST   : out    vl_logic;
        S09_AXI_RVALID  : out    vl_logic;
        S09_AXI_RREADY  : in     vl_logic;
        S10_AXI_ARESET_OUT_N: out    vl_logic;
        S10_AXI_ACLK    : in     vl_logic;
        S10_AXI_AWID    : in     vl_logic_vector;
        S10_AXI_AWADDR  : in     vl_logic_vector;
        S10_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S10_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S10_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S10_AXI_AWLOCK  : in     vl_logic;
        S10_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S10_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S10_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S10_AXI_AWVALID : in     vl_logic;
        S10_AXI_AWREADY : out    vl_logic;
        S10_AXI_WDATA   : in     vl_logic_vector;
        S10_AXI_WSTRB   : in     vl_logic_vector;
        S10_AXI_WLAST   : in     vl_logic;
        S10_AXI_WVALID  : in     vl_logic;
        S10_AXI_WREADY  : out    vl_logic;
        S10_AXI_BID     : out    vl_logic_vector;
        S10_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S10_AXI_BVALID  : out    vl_logic;
        S10_AXI_BREADY  : in     vl_logic;
        S10_AXI_ARID    : in     vl_logic_vector;
        S10_AXI_ARADDR  : in     vl_logic_vector;
        S10_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S10_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S10_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S10_AXI_ARLOCK  : in     vl_logic;
        S10_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S10_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S10_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S10_AXI_ARVALID : in     vl_logic;
        S10_AXI_ARREADY : out    vl_logic;
        S10_AXI_RID     : out    vl_logic_vector;
        S10_AXI_RDATA   : out    vl_logic_vector;
        S10_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S10_AXI_RLAST   : out    vl_logic;
        S10_AXI_RVALID  : out    vl_logic;
        S10_AXI_RREADY  : in     vl_logic;
        S11_AXI_ARESET_OUT_N: out    vl_logic;
        S11_AXI_ACLK    : in     vl_logic;
        S11_AXI_AWID    : in     vl_logic_vector;
        S11_AXI_AWADDR  : in     vl_logic_vector;
        S11_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S11_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S11_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S11_AXI_AWLOCK  : in     vl_logic;
        S11_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S11_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S11_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S11_AXI_AWVALID : in     vl_logic;
        S11_AXI_AWREADY : out    vl_logic;
        S11_AXI_WDATA   : in     vl_logic_vector;
        S11_AXI_WSTRB   : in     vl_logic_vector;
        S11_AXI_WLAST   : in     vl_logic;
        S11_AXI_WVALID  : in     vl_logic;
        S11_AXI_WREADY  : out    vl_logic;
        S11_AXI_BID     : out    vl_logic_vector;
        S11_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S11_AXI_BVALID  : out    vl_logic;
        S11_AXI_BREADY  : in     vl_logic;
        S11_AXI_ARID    : in     vl_logic_vector;
        S11_AXI_ARADDR  : in     vl_logic_vector;
        S11_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S11_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S11_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S11_AXI_ARLOCK  : in     vl_logic;
        S11_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S11_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S11_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S11_AXI_ARVALID : in     vl_logic;
        S11_AXI_ARREADY : out    vl_logic;
        S11_AXI_RID     : out    vl_logic_vector;
        S11_AXI_RDATA   : out    vl_logic_vector;
        S11_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S11_AXI_RLAST   : out    vl_logic;
        S11_AXI_RVALID  : out    vl_logic;
        S11_AXI_RREADY  : in     vl_logic;
        S12_AXI_ARESET_OUT_N: out    vl_logic;
        S12_AXI_ACLK    : in     vl_logic;
        S12_AXI_AWID    : in     vl_logic_vector;
        S12_AXI_AWADDR  : in     vl_logic_vector;
        S12_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S12_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S12_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S12_AXI_AWLOCK  : in     vl_logic;
        S12_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S12_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S12_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S12_AXI_AWVALID : in     vl_logic;
        S12_AXI_AWREADY : out    vl_logic;
        S12_AXI_WDATA   : in     vl_logic_vector;
        S12_AXI_WSTRB   : in     vl_logic_vector;
        S12_AXI_WLAST   : in     vl_logic;
        S12_AXI_WVALID  : in     vl_logic;
        S12_AXI_WREADY  : out    vl_logic;
        S12_AXI_BID     : out    vl_logic_vector;
        S12_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S12_AXI_BVALID  : out    vl_logic;
        S12_AXI_BREADY  : in     vl_logic;
        S12_AXI_ARID    : in     vl_logic_vector;
        S12_AXI_ARADDR  : in     vl_logic_vector;
        S12_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S12_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S12_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S12_AXI_ARLOCK  : in     vl_logic;
        S12_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S12_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S12_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S12_AXI_ARVALID : in     vl_logic;
        S12_AXI_ARREADY : out    vl_logic;
        S12_AXI_RID     : out    vl_logic_vector;
        S12_AXI_RDATA   : out    vl_logic_vector;
        S12_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S12_AXI_RLAST   : out    vl_logic;
        S12_AXI_RVALID  : out    vl_logic;
        S12_AXI_RREADY  : in     vl_logic;
        S13_AXI_ARESET_OUT_N: out    vl_logic;
        S13_AXI_ACLK    : in     vl_logic;
        S13_AXI_AWID    : in     vl_logic_vector;
        S13_AXI_AWADDR  : in     vl_logic_vector;
        S13_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S13_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S13_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S13_AXI_AWLOCK  : in     vl_logic;
        S13_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S13_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S13_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S13_AXI_AWVALID : in     vl_logic;
        S13_AXI_AWREADY : out    vl_logic;
        S13_AXI_WDATA   : in     vl_logic_vector;
        S13_AXI_WSTRB   : in     vl_logic_vector;
        S13_AXI_WLAST   : in     vl_logic;
        S13_AXI_WVALID  : in     vl_logic;
        S13_AXI_WREADY  : out    vl_logic;
        S13_AXI_BID     : out    vl_logic_vector;
        S13_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S13_AXI_BVALID  : out    vl_logic;
        S13_AXI_BREADY  : in     vl_logic;
        S13_AXI_ARID    : in     vl_logic_vector;
        S13_AXI_ARADDR  : in     vl_logic_vector;
        S13_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S13_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S13_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S13_AXI_ARLOCK  : in     vl_logic;
        S13_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S13_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S13_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S13_AXI_ARVALID : in     vl_logic;
        S13_AXI_ARREADY : out    vl_logic;
        S13_AXI_RID     : out    vl_logic_vector;
        S13_AXI_RDATA   : out    vl_logic_vector;
        S13_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S13_AXI_RLAST   : out    vl_logic;
        S13_AXI_RVALID  : out    vl_logic;
        S13_AXI_RREADY  : in     vl_logic;
        S14_AXI_ARESET_OUT_N: out    vl_logic;
        S14_AXI_ACLK    : in     vl_logic;
        S14_AXI_AWID    : in     vl_logic_vector;
        S14_AXI_AWADDR  : in     vl_logic_vector;
        S14_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S14_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S14_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S14_AXI_AWLOCK  : in     vl_logic;
        S14_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S14_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S14_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S14_AXI_AWVALID : in     vl_logic;
        S14_AXI_AWREADY : out    vl_logic;
        S14_AXI_WDATA   : in     vl_logic_vector;
        S14_AXI_WSTRB   : in     vl_logic_vector;
        S14_AXI_WLAST   : in     vl_logic;
        S14_AXI_WVALID  : in     vl_logic;
        S14_AXI_WREADY  : out    vl_logic;
        S14_AXI_BID     : out    vl_logic_vector;
        S14_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S14_AXI_BVALID  : out    vl_logic;
        S14_AXI_BREADY  : in     vl_logic;
        S14_AXI_ARID    : in     vl_logic_vector;
        S14_AXI_ARADDR  : in     vl_logic_vector;
        S14_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S14_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S14_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S14_AXI_ARLOCK  : in     vl_logic;
        S14_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S14_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S14_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S14_AXI_ARVALID : in     vl_logic;
        S14_AXI_ARREADY : out    vl_logic;
        S14_AXI_RID     : out    vl_logic_vector;
        S14_AXI_RDATA   : out    vl_logic_vector;
        S14_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S14_AXI_RLAST   : out    vl_logic;
        S14_AXI_RVALID  : out    vl_logic;
        S14_AXI_RREADY  : in     vl_logic;
        S15_AXI_ARESET_OUT_N: out    vl_logic;
        S15_AXI_ACLK    : in     vl_logic;
        S15_AXI_AWID    : in     vl_logic_vector;
        S15_AXI_AWADDR  : in     vl_logic_vector;
        S15_AXI_AWLEN   : in     vl_logic_vector(7 downto 0);
        S15_AXI_AWSIZE  : in     vl_logic_vector(2 downto 0);
        S15_AXI_AWBURST : in     vl_logic_vector(1 downto 0);
        S15_AXI_AWLOCK  : in     vl_logic;
        S15_AXI_AWCACHE : in     vl_logic_vector(3 downto 0);
        S15_AXI_AWPROT  : in     vl_logic_vector(2 downto 0);
        S15_AXI_AWQOS   : in     vl_logic_vector(3 downto 0);
        S15_AXI_AWVALID : in     vl_logic;
        S15_AXI_AWREADY : out    vl_logic;
        S15_AXI_WDATA   : in     vl_logic_vector;
        S15_AXI_WSTRB   : in     vl_logic_vector;
        S15_AXI_WLAST   : in     vl_logic;
        S15_AXI_WVALID  : in     vl_logic;
        S15_AXI_WREADY  : out    vl_logic;
        S15_AXI_BID     : out    vl_logic_vector;
        S15_AXI_BRESP   : out    vl_logic_vector(1 downto 0);
        S15_AXI_BVALID  : out    vl_logic;
        S15_AXI_BREADY  : in     vl_logic;
        S15_AXI_ARID    : in     vl_logic_vector;
        S15_AXI_ARADDR  : in     vl_logic_vector;
        S15_AXI_ARLEN   : in     vl_logic_vector(7 downto 0);
        S15_AXI_ARSIZE  : in     vl_logic_vector(2 downto 0);
        S15_AXI_ARBURST : in     vl_logic_vector(1 downto 0);
        S15_AXI_ARLOCK  : in     vl_logic;
        S15_AXI_ARCACHE : in     vl_logic_vector(3 downto 0);
        S15_AXI_ARPROT  : in     vl_logic_vector(2 downto 0);
        S15_AXI_ARQOS   : in     vl_logic_vector(3 downto 0);
        S15_AXI_ARVALID : in     vl_logic;
        S15_AXI_ARREADY : out    vl_logic;
        S15_AXI_RID     : out    vl_logic_vector;
        S15_AXI_RDATA   : out    vl_logic_vector;
        S15_AXI_RRESP   : out    vl_logic_vector(1 downto 0);
        S15_AXI_RLAST   : out    vl_logic;
        S15_AXI_RVALID  : out    vl_logic;
        S15_AXI_RREADY  : in     vl_logic;
        M00_AXI_ARESET_OUT_N: out    vl_logic;
        M00_AXI_ACLK    : in     vl_logic;
        M00_AXI_AWID    : out    vl_logic_vector;
        M00_AXI_AWADDR  : out    vl_logic_vector;
        M00_AXI_AWLEN   : out    vl_logic_vector(7 downto 0);
        M00_AXI_AWSIZE  : out    vl_logic_vector(2 downto 0);
        M00_AXI_AWBURST : out    vl_logic_vector(1 downto 0);
        M00_AXI_AWLOCK  : out    vl_logic;
        M00_AXI_AWCACHE : out    vl_logic_vector(3 downto 0);
        M00_AXI_AWPROT  : out    vl_logic_vector(2 downto 0);
        M00_AXI_AWQOS   : out    vl_logic_vector(3 downto 0);
        M00_AXI_AWVALID : out    vl_logic;
        M00_AXI_AWREADY : in     vl_logic;
        M00_AXI_WDATA   : out    vl_logic_vector;
        M00_AXI_WSTRB   : out    vl_logic_vector;
        M00_AXI_WLAST   : out    vl_logic;
        M00_AXI_WVALID  : out    vl_logic;
        M00_AXI_WREADY  : in     vl_logic;
        M00_AXI_BID     : in     vl_logic_vector;
        M00_AXI_BRESP   : in     vl_logic_vector(1 downto 0);
        M00_AXI_BVALID  : in     vl_logic;
        M00_AXI_BREADY  : out    vl_logic;
        M00_AXI_ARID    : out    vl_logic_vector;
        M00_AXI_ARADDR  : out    vl_logic_vector;
        M00_AXI_ARLEN   : out    vl_logic_vector(7 downto 0);
        M00_AXI_ARSIZE  : out    vl_logic_vector(2 downto 0);
        M00_AXI_ARBURST : out    vl_logic_vector(1 downto 0);
        M00_AXI_ARLOCK  : out    vl_logic;
        M00_AXI_ARCACHE : out    vl_logic_vector(3 downto 0);
        M00_AXI_ARPROT  : out    vl_logic_vector(2 downto 0);
        M00_AXI_ARQOS   : out    vl_logic_vector(3 downto 0);
        M00_AXI_ARVALID : out    vl_logic;
        M00_AXI_ARREADY : in     vl_logic;
        M00_AXI_RID     : in     vl_logic_vector;
        M00_AXI_RDATA   : in     vl_logic_vector;
        M00_AXI_RRESP   : in     vl_logic_vector(1 downto 0);
        M00_AXI_RLAST   : in     vl_logic;
        M00_AXI_RVALID  : in     vl_logic;
        M00_AXI_RREADY  : out    vl_logic
    );
end axi_interconnect_v1_06_a;
