library verilog;
use verilog.vl_types.all;
entity altpcietb_bfm_rp_top_x8_pipen1b is
    generic(
        RP_PRI_BUS_NUM  : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RP_PRI_DEV_NUM  : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        SHMEM_ADDR_WIDTH: integer := 21;
        EBFM_BAR_M64_MIN: vl_logic_vector(63 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EBFM_NUM_VC     : integer := 4;
        EBFM_NUM_TAG    : integer := 32;
        EBFM_MSG_DEBUG  : integer := 0;
        EBFM_MSG_INFO   : integer := 1;
        EBFM_MSG_WARNING: integer := 2;
        EBFM_MSG_ERROR_INFO: integer := 3;
        EBFM_MSG_ERROR_CONTINUE: integer := 4;
        EBFM_MSG_ERROR_FATAL: integer := 101;
        EBFM_MSG_ERROR_FATAL_TB_ERR: integer := 102;
        EBFM_MSG_MAX_LEN: integer := 100;
        SHMEM_FILL_ZERO : integer := 0;
        SHMEM_FILL_BYTE_INC: integer := 1;
        SHMEM_FILL_WORD_INC: integer := 2;
        SHMEM_FILL_DWORD_INC: integer := 4;
        SHMEM_FILL_QWORD_INC: integer := 8;
        SHMEM_FILL_ONE  : integer := 15;
        BAR_TABLE_SIZE  : integer := 64;
        SCR_SIZE        : integer := 64
    );
    port(
        clk250_in       : in     vl_logic;
        clk500_in       : in     vl_logic;
        local_rstn      : in     vl_logic;
        pcie_rstn       : in     vl_logic;
        swdn_out        : out    vl_logic_vector(5 downto 0);
        rx_in0          : in     vl_logic;
        tx_out0         : out    vl_logic;
        rx_in1          : in     vl_logic;
        tx_out1         : out    vl_logic;
        rx_in2          : in     vl_logic;
        tx_out2         : out    vl_logic;
        rx_in3          : in     vl_logic;
        tx_out3         : out    vl_logic;
        rx_in4          : in     vl_logic;
        tx_out4         : out    vl_logic;
        rx_in5          : in     vl_logic;
        tx_out5         : out    vl_logic;
        rx_in6          : in     vl_logic;
        tx_out6         : out    vl_logic;
        rx_in7          : in     vl_logic;
        tx_out7         : out    vl_logic;
        pipe_mode       : in     vl_logic;
        test_in         : in     vl_logic_vector(31 downto 0);
        test_out        : out    vl_logic_vector(511 downto 0);
        txdata0_ext     : out    vl_logic_vector(7 downto 0);
        txdatak0_ext    : out    vl_logic;
        txdetectrx0_ext : out    vl_logic;
        txelecidle0_ext : out    vl_logic;
        txcompl0_ext    : out    vl_logic;
        rxpolarity0_ext : out    vl_logic;
        powerdown0_ext  : out    vl_logic_vector(1 downto 0);
        rxdata0_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak0_ext    : in     vl_logic;
        rxvalid0_ext    : in     vl_logic;
        phystatus0_ext  : in     vl_logic;
        rxelecidle0_ext : in     vl_logic;
        rxstatus0_ext   : in     vl_logic_vector(2 downto 0);
        txdata1_ext     : out    vl_logic_vector(7 downto 0);
        txdatak1_ext    : out    vl_logic;
        txdetectrx1_ext : out    vl_logic;
        txelecidle1_ext : out    vl_logic;
        txcompl1_ext    : out    vl_logic;
        rxpolarity1_ext : out    vl_logic;
        powerdown1_ext  : out    vl_logic_vector(1 downto 0);
        rxdata1_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak1_ext    : in     vl_logic;
        rxvalid1_ext    : in     vl_logic;
        phystatus1_ext  : in     vl_logic;
        rxelecidle1_ext : in     vl_logic;
        rxstatus1_ext   : in     vl_logic_vector(2 downto 0);
        txdata2_ext     : out    vl_logic_vector(7 downto 0);
        txdatak2_ext    : out    vl_logic;
        txdetectrx2_ext : out    vl_logic;
        txelecidle2_ext : out    vl_logic;
        txcompl2_ext    : out    vl_logic;
        rxpolarity2_ext : out    vl_logic;
        powerdown2_ext  : out    vl_logic_vector(1 downto 0);
        rxdata2_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak2_ext    : in     vl_logic;
        rxvalid2_ext    : in     vl_logic;
        phystatus2_ext  : in     vl_logic;
        rxelecidle2_ext : in     vl_logic;
        rxstatus2_ext   : in     vl_logic_vector(2 downto 0);
        txdata3_ext     : out    vl_logic_vector(7 downto 0);
        txdatak3_ext    : out    vl_logic;
        txdetectrx3_ext : out    vl_logic;
        txelecidle3_ext : out    vl_logic;
        txcompl3_ext    : out    vl_logic;
        rxpolarity3_ext : out    vl_logic;
        powerdown3_ext  : out    vl_logic_vector(1 downto 0);
        rxdata3_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak3_ext    : in     vl_logic;
        rxvalid3_ext    : in     vl_logic;
        phystatus3_ext  : in     vl_logic;
        rxelecidle3_ext : in     vl_logic;
        rxstatus3_ext   : in     vl_logic_vector(2 downto 0);
        txdata4_ext     : out    vl_logic_vector(7 downto 0);
        txdatak4_ext    : out    vl_logic;
        txdetectrx4_ext : out    vl_logic;
        txelecidle4_ext : out    vl_logic;
        txcompl4_ext    : out    vl_logic;
        rxpolarity4_ext : out    vl_logic;
        powerdown4_ext  : out    vl_logic_vector(1 downto 0);
        rxdata4_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak4_ext    : in     vl_logic;
        rxvalid4_ext    : in     vl_logic;
        phystatus4_ext  : in     vl_logic;
        rxelecidle4_ext : in     vl_logic;
        rxstatus4_ext   : in     vl_logic_vector(2 downto 0);
        txdata5_ext     : out    vl_logic_vector(7 downto 0);
        txdatak5_ext    : out    vl_logic;
        txdetectrx5_ext : out    vl_logic;
        txelecidle5_ext : out    vl_logic;
        txcompl5_ext    : out    vl_logic;
        rxpolarity5_ext : out    vl_logic;
        powerdown5_ext  : out    vl_logic_vector(1 downto 0);
        rxdata5_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak5_ext    : in     vl_logic;
        rxvalid5_ext    : in     vl_logic;
        phystatus5_ext  : in     vl_logic;
        rxelecidle5_ext : in     vl_logic;
        rxstatus5_ext   : in     vl_logic_vector(2 downto 0);
        txdata6_ext     : out    vl_logic_vector(7 downto 0);
        txdatak6_ext    : out    vl_logic;
        txdetectrx6_ext : out    vl_logic;
        txelecidle6_ext : out    vl_logic;
        txcompl6_ext    : out    vl_logic;
        rxpolarity6_ext : out    vl_logic;
        powerdown6_ext  : out    vl_logic_vector(1 downto 0);
        rxdata6_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak6_ext    : in     vl_logic;
        rxvalid6_ext    : in     vl_logic;
        phystatus6_ext  : in     vl_logic;
        rxelecidle6_ext : in     vl_logic;
        rxstatus6_ext   : in     vl_logic_vector(2 downto 0);
        txdata7_ext     : out    vl_logic_vector(7 downto 0);
        txdatak7_ext    : out    vl_logic;
        txdetectrx7_ext : out    vl_logic;
        txelecidle7_ext : out    vl_logic;
        txcompl7_ext    : out    vl_logic;
        rxpolarity7_ext : out    vl_logic;
        powerdown7_ext  : out    vl_logic_vector(1 downto 0);
        rxdata7_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak7_ext    : in     vl_logic;
        rxvalid7_ext    : in     vl_logic;
        phystatus7_ext  : in     vl_logic;
        rxelecidle7_ext : in     vl_logic;
        rxstatus7_ext   : in     vl_logic_vector(2 downto 0);
        rate_ext        : out    vl_logic
    );
    attribute RP_PRI_BUS_NUM_mti_vect_attrib : integer;
    attribute RP_PRI_BUS_NUM_mti_vect_attrib of RP_PRI_BUS_NUM : constant is 0;
    attribute RP_PRI_DEV_NUM_mti_vect_attrib : integer;
    attribute RP_PRI_DEV_NUM_mti_vect_attrib of RP_PRI_DEV_NUM : constant is 0;
    attribute EBFM_BAR_M64_MIN_mti_vect_attrib : integer;
    attribute EBFM_BAR_M64_MIN_mti_vect_attrib of EBFM_BAR_M64_MIN : constant is 0;
end altpcietb_bfm_rp_top_x8_pipen1b;
