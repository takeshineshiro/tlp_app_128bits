library verilog;
use verilog.vl_types.all;
entity ict106_converter_bank is
    generic(
        C_FAMILY        : string  := "none";
        C_NUM_SLOTS     : integer := 1;
        C_AXI_ID_WIDTH  : integer := 1;
        C_AXI_ID_MAX_WIDTH: integer := 1;
        C_AXI_ADDR_WIDTH: integer := 32;
        C_AXI_DATA_MAX_WIDTH: integer := 256;
        C_AXI_PROTOCOL  : integer := 0;
        C_AXI_IS_ACLK_ASYNC: integer := 0;
        C_AXI_SUPPORTS_WRITE: integer := 65535;
        C_AXI_SUPPORTS_READ: integer := 65535;
        C_AXI_SUPPORTS_USER_SIGNALS: integer := 0;
        C_AXI_AWUSER_WIDTH: integer := 1;
        C_AXI_ARUSER_WIDTH: integer := 1;
        C_AXI_WUSER_WIDTH: integer := 1;
        C_AXI_RUSER_WIDTH: integer := 1;
        C_AXI_BUSER_WIDTH: integer := 1;
        C_HEMISPHERE    : string  := "si"
    );
    port(
        INTERCONNECT_ACLK: in     vl_logic;
        INTERCONNECT_ARESETN: in     vl_logic;
        LOCAL_ARESETN   : in     vl_logic;
        INTERCONNECT_RESET_OUT_N: out    vl_logic;
        S_AXI_RESET_OUT_N: out    vl_logic_vector;
        M_AXI_RESET_OUT_N: out    vl_logic_vector;
        S_AXI_ACLK      : in     vl_logic_vector;
        S_AXI_AWID      : in     vl_logic_vector;
        S_AXI_AWADDR    : in     vl_logic_vector;
        S_AXI_AWLEN     : in     vl_logic_vector;
        S_AXI_AWSIZE    : in     vl_logic_vector;
        S_AXI_AWBURST   : in     vl_logic_vector;
        S_AXI_AWLOCK    : in     vl_logic_vector;
        S_AXI_AWCACHE   : in     vl_logic_vector;
        S_AXI_AWPROT    : in     vl_logic_vector;
        S_AXI_AWREGION  : in     vl_logic_vector;
        S_AXI_AWQOS     : in     vl_logic_vector;
        S_AXI_AWUSER    : in     vl_logic_vector;
        S_AXI_AWVALID   : in     vl_logic_vector;
        S_AXI_AWREADY   : out    vl_logic_vector;
        S_AXI_WDATA     : in     vl_logic_vector;
        S_AXI_WSTRB     : in     vl_logic_vector;
        S_AXI_WLAST     : in     vl_logic_vector;
        S_AXI_WUSER     : in     vl_logic_vector;
        S_AXI_WVALID    : in     vl_logic_vector;
        S_AXI_WREADY    : out    vl_logic_vector;
        S_AXI_BID       : out    vl_logic_vector;
        S_AXI_BRESP     : out    vl_logic_vector;
        S_AXI_BUSER     : out    vl_logic_vector;
        S_AXI_BVALID    : out    vl_logic_vector;
        S_AXI_BREADY    : in     vl_logic_vector;
        S_AXI_ARID      : in     vl_logic_vector;
        S_AXI_ARADDR    : in     vl_logic_vector;
        S_AXI_ARLEN     : in     vl_logic_vector;
        S_AXI_ARSIZE    : in     vl_logic_vector;
        S_AXI_ARBURST   : in     vl_logic_vector;
        S_AXI_ARLOCK    : in     vl_logic_vector;
        S_AXI_ARCACHE   : in     vl_logic_vector;
        S_AXI_ARPROT    : in     vl_logic_vector;
        S_AXI_ARREGION  : in     vl_logic_vector;
        S_AXI_ARQOS     : in     vl_logic_vector;
        S_AXI_ARUSER    : in     vl_logic_vector;
        S_AXI_ARVALID   : in     vl_logic_vector;
        S_AXI_ARREADY   : out    vl_logic_vector;
        S_AXI_RID       : out    vl_logic_vector;
        S_AXI_RDATA     : out    vl_logic_vector;
        S_AXI_RRESP     : out    vl_logic_vector;
        S_AXI_RLAST     : out    vl_logic_vector;
        S_AXI_RUSER     : out    vl_logic_vector;
        S_AXI_RVALID    : out    vl_logic_vector;
        S_AXI_RREADY    : in     vl_logic_vector;
        M_AXI_ACLK      : in     vl_logic_vector;
        M_AXI_AWID      : out    vl_logic_vector;
        M_AXI_AWADDR    : out    vl_logic_vector;
        M_AXI_AWLEN     : out    vl_logic_vector;
        M_AXI_AWSIZE    : out    vl_logic_vector;
        M_AXI_AWBURST   : out    vl_logic_vector;
        M_AXI_AWLOCK    : out    vl_logic_vector;
        M_AXI_AWCACHE   : out    vl_logic_vector;
        M_AXI_AWPROT    : out    vl_logic_vector;
        M_AXI_AWREGION  : out    vl_logic_vector;
        M_AXI_AWQOS     : out    vl_logic_vector;
        M_AXI_AWUSER    : out    vl_logic_vector;
        M_AXI_AWVALID   : out    vl_logic_vector;
        M_AXI_AWREADY   : in     vl_logic_vector;
        M_AXI_WDATA     : out    vl_logic_vector;
        M_AXI_WSTRB     : out    vl_logic_vector;
        M_AXI_WLAST     : out    vl_logic_vector;
        M_AXI_WUSER     : out    vl_logic_vector;
        M_AXI_WVALID    : out    vl_logic_vector;
        M_AXI_WREADY    : in     vl_logic_vector;
        M_AXI_BID       : in     vl_logic_vector;
        M_AXI_BRESP     : in     vl_logic_vector;
        M_AXI_BUSER     : in     vl_logic_vector;
        M_AXI_BVALID    : in     vl_logic_vector;
        M_AXI_BREADY    : out    vl_logic_vector;
        M_AXI_ARID      : out    vl_logic_vector;
        M_AXI_ARADDR    : out    vl_logic_vector;
        M_AXI_ARLEN     : out    vl_logic_vector;
        M_AXI_ARSIZE    : out    vl_logic_vector;
        M_AXI_ARBURST   : out    vl_logic_vector;
        M_AXI_ARLOCK    : out    vl_logic_vector;
        M_AXI_ARCACHE   : out    vl_logic_vector;
        M_AXI_ARPROT    : out    vl_logic_vector;
        M_AXI_ARREGION  : out    vl_logic_vector;
        M_AXI_ARQOS     : out    vl_logic_vector;
        M_AXI_ARUSER    : out    vl_logic_vector;
        M_AXI_ARVALID   : out    vl_logic_vector;
        M_AXI_ARREADY   : in     vl_logic_vector;
        M_AXI_RID       : in     vl_logic_vector;
        M_AXI_RDATA     : in     vl_logic_vector;
        M_AXI_RRESP     : in     vl_logic_vector;
        M_AXI_RLAST     : in     vl_logic_vector;
        M_AXI_RUSER     : in     vl_logic_vector;
        M_AXI_RVALID    : in     vl_logic_vector;
        M_AXI_RREADY    : out    vl_logic_vector
    );
end ict106_converter_bank;
