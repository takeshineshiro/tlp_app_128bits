// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: scfifo 

// ============================================================
// File Name: fifo.v
// Megafunction Name(s):
// 			scfifo
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 173 11/01/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module fifo (
	aclr,
	clock,
	data,
	rdreq,
	sclr,
	wrreq,
	almost_empty,
	almost_full,
	empty,
	full,
	q,
	usedw);
   parameter MEM_TYPE = 1;
   parameter DATA_W = 32;
   parameter DEPTH_W = 9;
	input	  aclr;
	input	  clock;
	input	[DATA_W-1:0]  data;
	input	  rdreq;
	input	  sclr;
	input	  wrreq;
	output	  almost_empty;
	output	  almost_full;
	output	  empty;
	output	  full;
	output	[DATA_W-1:0]  q;
	output	[DEPTH_W-1:0]  usedw;

	wire [DEPTH_W-1:0] sub_wire0;
	wire  sub_wire1;
	wire  sub_wire2;
	wire [DATA_W-1:0] sub_wire3;
	wire  sub_wire4;
	wire  sub_wire5;
	wire [DEPTH_W-1:0] usedw = sub_wire0[DEPTH_W-1:0];
	wire  empty = sub_wire1;
	wire  full = sub_wire2;
	wire [DATA_W-1:0] q = sub_wire3[DATA_W-1:0];
	wire  almost_empty = sub_wire4;
	wire  almost_full = sub_wire5;

	scfifo	scfifo_component (
				.clock (clock),
				.sclr (sclr),
				.wrreq (wrreq),
				.aclr (aclr),
				.data (data),
				.rdreq (rdreq),
				.usedw (sub_wire0),
				.empty (sub_wire1),
				.full (sub_wire2),
				.q (sub_wire3),
				.almost_empty (sub_wire4),
				.almost_full (sub_wire5));

	defparam
		scfifo_component.add_ram_output_register = "OFF",
		scfifo_component.almost_empty_value = 1,
		scfifo_component.almost_full_value = 1,
		scfifo_component.intended_device_family = "Stratix IV",
		scfifo_component.lpm_numwords = (1 << DEPTH_W),
		scfifo_component.lpm_showahead = "ON",
		scfifo_component.lpm_type = "scfifo",
		scfifo_component.lpm_width = DATA_W,
		scfifo_component.lpm_widthu = DEPTH_W,
		scfifo_component.overflow_checking = "ON",
		scfifo_component.underflow_checking = "ON",
		scfifo_component.use_eab = "ON";

endmodule



