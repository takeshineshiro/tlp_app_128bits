library verilog;
use verilog.vl_types.all;
entity axi_pcie is
    generic(
        C_INSTANCE      : string  := "AXI_PCIe";
        C_MAX_LINK_SPEED: integer := 0;
        C_PCIE_USE_MODE : string  := "1.0";
        C_DEVICE_ID     : integer := 4;
        C_VENDOR_ID     : integer := 4466;
        C_REV_ID        : integer := 1;
        C_SUBSYSTEM_ID  : integer := 0;
        C_SUBSYSTEM_VENDOR_ID: integer := 0;
        C_CLASS_CODE    : integer := 0;
        C_REF_CLK_FREQ  : integer := 0;
        C_PCIE_CAP_SLOT_IMPLEMENTED: integer := 0;
        C_NUM_MSI_REQ   : integer := 0;
        C_INTERRUPT_PIN : integer := 0;
        C_BASEADDR      : integer := -1;
        C_HIGHADDR      : integer := 0;
        C_NO_OF_LANES   : integer := 4;
        C_FAMILY        : string  := "virtex6";
        C_S_AXI_ID_WIDTH: integer := 4;
        C_S_AXI_ADDR_WIDTH: integer := 32;
        C_S_AXI_DATA_WIDTH: integer := 32;
        C_M_AXI_ADDR_WIDTH: integer := 32;
        C_M_AXI_DATA_WIDTH: integer := 32;
        C_COMP_TIMEOUT  : integer := 0;
        C_INCLUDE_RC    : integer := 0;
        C_S_AXI_SUPPORTS_NARROW_BURST: integer := 1;
        C_INCLUDE_BAROFFSET_REG: integer := 1;
        C_AXIBAR_NUM    : integer := 6;
        C_AXIBAR2PCIEBAR_0: integer := 0;
        C_AXIBAR2PCIEBAR_1: integer := 0;
        C_AXIBAR2PCIEBAR_2: integer := 0;
        C_AXIBAR2PCIEBAR_3: integer := 0;
        C_AXIBAR2PCIEBAR_4: integer := 0;
        C_AXIBAR2PCIEBAR_5: integer := 0;
        C_AXIBAR_AS_0   : integer := 0;
        C_AXIBAR_AS_1   : integer := 0;
        C_AXIBAR_AS_2   : integer := 0;
        C_AXIBAR_AS_3   : integer := 0;
        C_AXIBAR_AS_4   : integer := 0;
        C_AXIBAR_AS_5   : integer := 0;
        C_AXIBAR_0      : integer := -1;
        C_AXIBAR_HIGHADDR_0: integer := 0;
        C_AXIBAR_1      : integer := -1;
        C_AXIBAR_HIGHADDR_1: integer := 0;
        C_AXIBAR_2      : integer := -1;
        C_AXIBAR_HIGHADDR_2: integer := 0;
        C_AXIBAR_3      : integer := -1;
        C_AXIBAR_HIGHADDR_3: integer := 0;
        C_AXIBAR_4      : integer := -1;
        C_AXIBAR_HIGHADDR_4: integer := 0;
        C_AXIBAR_5      : integer := -1;
        C_AXIBAR_HIGHADDR_5: integer := 0;
        C_PCIEBAR_NUM   : integer := 3;
        C_PCIEBAR_AS    : integer := 1;
        C_PCIEBAR_LEN_0 : integer := 16;
        C_PCIEBAR2AXIBAR_0: integer := 0;
        C_PCIEBAR_LEN_1 : integer := 16;
        C_PCIEBAR2AXIBAR_1: integer := 0;
        C_PCIEBAR_LEN_2 : integer := 16;
        C_PCIEBAR2AXIBAR_2: integer := 0;
        C_PIPE_MODE     : integer := 0;
        PCIE_BRAM_DEBUG_EN: integer := 0
    );
    port(
        linkdown        : out    vl_logic;
        clk_50M_out     : out    vl_logic;
        pll_locked      : out    vl_logic;
        axi_aclk_out    : out    vl_logic;
        axi_aresetn_out : out    vl_logic;
        pci_exp_txp     : out    vl_logic_vector;
        pci_exp_txn     : out    vl_logic_vector;
        axi_ctl_aclk_out: out    vl_logic;
        mmcm_lock       : out    vl_logic;
        interrupt_out   : out    vl_logic;
        INTX_MSI_Grant  : out    vl_logic;
        MSI_enable      : out    vl_logic;
        MSI_Vector_Width: out    vl_logic;
        s_axi_ctl_awready: out    vl_logic;
        s_axi_ctl_wready: out    vl_logic;
        s_axi_ctl_bresp : out    vl_logic_vector(1 downto 0);
        s_axi_ctl_bvalid: out    vl_logic;
        s_axi_ctl_arready: out    vl_logic;
        s_axi_ctl_rdata : out    vl_logic_vector(31 downto 0);
        s_axi_ctl_rresp : out    vl_logic_vector(1 downto 0);
        s_axi_ctl_rvalid: out    vl_logic;
        s_axi_awready   : out    vl_logic;
        s_axi_wready    : out    vl_logic;
        s_axi_bid       : out    vl_logic_vector;
        s_axi_bresp     : out    vl_logic_vector(1 downto 0);
        s_axi_bvalid    : out    vl_logic;
        s_axi_arready   : out    vl_logic;
        s_axi_rdata     : out    vl_logic_vector;
        s_axi_rid       : out    vl_logic_vector;
        s_axi_rresp     : out    vl_logic_vector(1 downto 0);
        s_axi_rlast     : out    vl_logic;
        s_axi_rvalid    : out    vl_logic;
        m_axi_awaddr    : out    vl_logic_vector;
        m_axi_awregion  : out    vl_logic_vector(3 downto 0);
        m_axi_awlen     : out    vl_logic_vector(7 downto 0);
        m_axi_awsize    : out    vl_logic_vector(2 downto 0);
        m_axi_awburst   : out    vl_logic_vector(1 downto 0);
        m_axi_awvalid   : out    vl_logic;
        m_axi_awcache   : out    vl_logic_vector(3 downto 0);
        m_axi_awlock    : out    vl_logic;
        m_axi_awprot    : out    vl_logic_vector(2 downto 0);
        m_axi_arlock    : out    vl_logic;
        m_axi_arcache   : out    vl_logic_vector(3 downto 0);
        m_axi_wdata     : out    vl_logic_vector;
        m_axi_wstrb     : out    vl_logic_vector;
        m_axi_wlast     : out    vl_logic;
        m_axi_wvalid    : out    vl_logic;
        m_axi_bready    : out    vl_logic;
        m_axi_arid      : out    vl_logic_vector;
        m_axi_araddr    : out    vl_logic_vector;
        m_axi_arregion  : out    vl_logic_vector(3 downto 0);
        m_axi_arlen     : out    vl_logic_vector(7 downto 0);
        m_axi_arsize    : out    vl_logic_vector(2 downto 0);
        m_axi_arburst   : out    vl_logic_vector(1 downto 0);
        m_axi_arvalid   : out    vl_logic;
        m_axi_arprot    : out    vl_logic_vector(2 downto 0);
        m_axi_rready    : out    vl_logic;
        m_axi_awready_user: out    vl_logic;
        m_axi_wready_user: out    vl_logic;
        m_axi_bresp_user: out    vl_logic_vector(1 downto 0);
        m_axi_bvalid_user: out    vl_logic;
        m_axi_arready_user: out    vl_logic;
        m_axi_rdata_user: out    vl_logic_vector(31 downto 0);
        m_axi_rresp_user: out    vl_logic_vector(1 downto 0);
        m_axi_rvalid_user: out    vl_logic;
        core_clk_out    : out    vl_logic;
        app_rst         : out    vl_logic;
        test_out_icm    : out    vl_logic_vector(8 downto 0);
        powerdown_ext   : out    vl_logic_vector(1 downto 0);
        rate_ext        : out    vl_logic;
        clk250_out      : out    vl_logic;
        clk500_out      : out    vl_logic;
        rxpolarity0_ext : out    vl_logic;
        txcompl0_ext    : out    vl_logic;
        txdata0_ext     : out    vl_logic_vector(7 downto 0);
        txdatak0_ext    : out    vl_logic;
        txelecidle0_ext : out    vl_logic;
        rxpolarity1_ext : out    vl_logic;
        txcompl1_ext    : out    vl_logic;
        txdata1_ext     : out    vl_logic_vector(7 downto 0);
        txdatak1_ext    : out    vl_logic;
        txelecidle1_ext : out    vl_logic;
        rxpolarity2_ext : out    vl_logic;
        txcompl2_ext    : out    vl_logic;
        txdata2_ext     : out    vl_logic_vector(7 downto 0);
        txdatak2_ext    : out    vl_logic;
        txelecidle2_ext : out    vl_logic;
        rxpolarity3_ext : out    vl_logic;
        txcompl3_ext    : out    vl_logic;
        txdata3_ext     : out    vl_logic_vector(7 downto 0);
        txdatak3_ext    : out    vl_logic;
        txelecidle3_ext : out    vl_logic;
        rxpolarity4_ext : out    vl_logic;
        txcompl4_ext    : out    vl_logic;
        txdata4_ext     : out    vl_logic_vector(7 downto 0);
        txdatak4_ext    : out    vl_logic;
        txelecidle4_ext : out    vl_logic;
        rxpolarity5_ext : out    vl_logic;
        txcompl5_ext    : out    vl_logic;
        txdata5_ext     : out    vl_logic_vector(7 downto 0);
        txdatak5_ext    : out    vl_logic;
        txelecidle5_ext : out    vl_logic;
        rxpolarity6_ext : out    vl_logic;
        txcompl6_ext    : out    vl_logic;
        txdata6_ext     : out    vl_logic_vector(7 downto 0);
        txdatak6_ext    : out    vl_logic;
        txelecidle6_ext : out    vl_logic;
        rxpolarity7_ext : out    vl_logic;
        txcompl7_ext    : out    vl_logic;
        txdata7_ext     : out    vl_logic_vector(7 downto 0);
        txdatak7_ext    : out    vl_logic;
        txelecidle7_ext : out    vl_logic;
        txdetectrx_ext  : out    vl_logic;
        free_100MHz     : in     vl_logic;
        pcie_rstn       : in     vl_logic;
        axi_aclk        : in     vl_logic;
        axi_aresetn     : in     vl_logic;
        INTX_MSI_Request: in     vl_logic;
        REFCLK          : in     vl_logic;
        pci_exp_rxp     : in     vl_logic_vector;
        pci_exp_rxn     : in     vl_logic_vector;
        axi_ctl_aclk    : in     vl_logic;
        MSI_Vector_Num  : in     vl_logic;
        s_axi_ctl_awaddr: in     vl_logic_vector(31 downto 0);
        s_axi_ctl_awvalid: in     vl_logic;
        s_axi_ctl_wdata : in     vl_logic_vector(31 downto 0);
        s_axi_ctl_wstrb : in     vl_logic_vector(3 downto 0);
        s_axi_ctl_wvalid: in     vl_logic;
        s_axi_ctl_bready: in     vl_logic;
        s_axi_ctl_araddr: in     vl_logic_vector(31 downto 0);
        s_axi_ctl_arvalid: in     vl_logic;
        s_axi_ctl_rready: in     vl_logic;
        s_axi_awid      : in     vl_logic_vector;
        s_axi_awaddr    : in     vl_logic_vector;
        s_axi_awregion  : in     vl_logic_vector(3 downto 0);
        s_axi_awlen     : in     vl_logic_vector(7 downto 0);
        s_axi_awsize    : in     vl_logic_vector(2 downto 0);
        s_axi_awburst   : in     vl_logic_vector(1 downto 0);
        s_axi_awvalid   : in     vl_logic;
        s_axi_wdata     : in     vl_logic_vector;
        s_axi_wstrb     : in     vl_logic_vector;
        s_axi_wlast     : in     vl_logic;
        s_axi_wvalid    : in     vl_logic;
        s_axi_bready    : in     vl_logic;
        s_axi_arid      : in     vl_logic_vector;
        s_axi_araddr    : in     vl_logic_vector;
        s_axi_arregion  : in     vl_logic_vector(3 downto 0);
        s_axi_arlen     : in     vl_logic_vector(7 downto 0);
        s_axi_arsize    : in     vl_logic_vector(2 downto 0);
        s_axi_arburst   : in     vl_logic_vector(1 downto 0);
        s_axi_arvalid   : in     vl_logic;
        s_axi_rready    : in     vl_logic;
        m_axi_awready   : in     vl_logic;
        m_axi_wready    : in     vl_logic;
        m_axi_bresp     : in     vl_logic_vector(1 downto 0);
        m_axi_bvalid    : in     vl_logic;
        m_axi_arready   : in     vl_logic;
        m_axi_rdata     : in     vl_logic_vector;
        m_axi_rid       : in     vl_logic_vector;
        m_axi_rresp     : in     vl_logic_vector(1 downto 0);
        m_axi_rlast     : in     vl_logic;
        m_axi_rvalid    : in     vl_logic;
        m_axi_awvalid_user: in     vl_logic;
        m_axi_awaddr_user: in     vl_logic_vector(31 downto 0);
        m_axi_wdata_user: in     vl_logic_vector(31 downto 0);
        m_axi_wvalid_user: in     vl_logic;
        m_axi_bready_user: in     vl_logic;
        m_axi_arvalid_user: in     vl_logic;
        m_axi_araddr_user: in     vl_logic_vector(31 downto 0);
        m_axi_rready_user: in     vl_logic;
        test_in         : in     vl_logic_vector(39 downto 0);
        phystatus_ext   : in     vl_logic;
        pclk_in         : in     vl_logic;
        rxdata0_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak0_ext    : in     vl_logic;
        rxelecidle0_ext : in     vl_logic;
        rxstatus0_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid0_ext    : in     vl_logic;
        rxdata1_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak1_ext    : in     vl_logic;
        rxelecidle1_ext : in     vl_logic;
        rxstatus1_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid1_ext    : in     vl_logic;
        rxdata2_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak2_ext    : in     vl_logic;
        rxelecidle2_ext : in     vl_logic;
        rxstatus2_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid2_ext    : in     vl_logic;
        rxdata3_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak3_ext    : in     vl_logic;
        rxelecidle3_ext : in     vl_logic;
        rxstatus3_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid3_ext    : in     vl_logic;
        rxdata4_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak4_ext    : in     vl_logic;
        rxelecidle4_ext : in     vl_logic;
        rxstatus4_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid4_ext    : in     vl_logic;
        rxdata5_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak5_ext    : in     vl_logic;
        rxelecidle5_ext : in     vl_logic;
        rxstatus5_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid5_ext    : in     vl_logic;
        rxdata6_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak6_ext    : in     vl_logic;
        rxelecidle6_ext : in     vl_logic;
        rxstatus6_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid6_ext    : in     vl_logic;
        rxdata7_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak7_ext    : in     vl_logic;
        rxelecidle7_ext : in     vl_logic;
        rxstatus7_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid7_ext    : in     vl_logic
    );
end axi_pcie;
