library verilog;
use verilog.vl_types.all;
entity pcie_top is
    generic(
        PCIE_VENDOR_ID  : integer := 4466;
        PCIE_DEVICE_ID  : integer := 4;
        PCIE_VEVISION_ID: integer := 1
    );
    port(
        pcie_rstn       : in     vl_logic;
        refclk          : in     vl_logic;
        app_rst         : out    vl_logic;
        core_clk_out    : out    vl_logic;
        rx_in0          : in     vl_logic;
        tx_out0         : out    vl_logic;
        rx_in1          : in     vl_logic;
        rx_in2          : in     vl_logic;
        rx_in3          : in     vl_logic;
        tx_out1         : out    vl_logic;
        tx_out2         : out    vl_logic;
        tx_out3         : out    vl_logic;
        rx_in4          : in     vl_logic;
        rx_in5          : in     vl_logic;
        rx_in6          : in     vl_logic;
        rx_in7          : in     vl_logic;
        tx_out4         : out    vl_logic;
        tx_out5         : out    vl_logic;
        tx_out6         : out    vl_logic;
        tx_out7         : out    vl_logic;
        app_int_ack     : out    vl_logic;
        app_int_sts     : in     vl_logic;
        app_msi_ack     : out    vl_logic;
        app_msi_num     : in     vl_logic_vector(4 downto 0);
        app_msi_req     : in     vl_logic;
        app_msi_tc      : in     vl_logic_vector(2 downto 0);
        pex_msi_num     : in     vl_logic_vector(4 downto 0);
        rx_fifo_empty0  : out    vl_logic;
        rx_fifo_full0   : out    vl_logic;
        rx_st_err0      : out    vl_logic;
        rx_st_bardec0   : out    vl_logic_vector(7 downto 0);
        rx_st_data0     : out    vl_logic_vector(63 downto 0);
        rx_st_be0       : out    vl_logic_vector(7 downto 0);
        rx_st_sop0      : out    vl_logic;
        rx_st_eop0      : out    vl_logic;
        rx_st_ready0    : in     vl_logic;
        rx_st_valid0    : out    vl_logic;
        tx_cred0        : out    vl_logic_vector(35 downto 0);
        tx_fifo_empty0  : out    vl_logic;
        tx_fifo_full0   : out    vl_logic;
        tx_fifo_rdptr0  : out    vl_logic_vector(3 downto 0);
        tx_fifo_wrptr0  : out    vl_logic_vector(3 downto 0);
        tx_st_data0     : in     vl_logic_vector(63 downto 0);
        tx_st_sop0      : in     vl_logic;
        tx_st_eop0      : in     vl_logic;
        tx_st_ready0    : out    vl_logic;
        tx_st_valid0    : in     vl_logic;
        linkdown        : out    vl_logic;
        gen2_led        : out    vl_logic;
        maxpayloadsize  : out    vl_logic_vector(2 downto 0);
        maxreadrequestsize: out    vl_logic_vector(2 downto 0);
        completerid     : out    vl_logic_vector(12 downto 0);
        cpl_pending     : in     vl_logic;
        cpl_err_in      : in     vl_logic_vector(6 downto 0);
        reconfig_clk_locked: in     vl_logic;
        reconfig_clk    : in     vl_logic;
        fixedclk_serdes : in     vl_logic;
        test_in         : in     vl_logic_vector(39 downto 0);
        test_out        : out    vl_logic_vector(8 downto 0);
        lane_act        : out    vl_logic_vector(3 downto 0);
        pipe_mode       : in     vl_logic;
        powerdown_ext   : out    vl_logic_vector(1 downto 0);
        phystatus_ext   : in     vl_logic;
        rate_ext        : out    vl_logic;
        pclk_in         : in     vl_logic;
        clk250_out      : out    vl_logic;
        clk500_out      : out    vl_logic;
        rxdata0_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak0_ext    : in     vl_logic;
        rxelecidle0_ext : in     vl_logic;
        rxpolarity0_ext : out    vl_logic;
        rxstatus0_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid0_ext    : in     vl_logic;
        txcompl0_ext    : out    vl_logic;
        txdata0_ext     : out    vl_logic_vector(7 downto 0);
        txdatak0_ext    : out    vl_logic;
        txelecidle0_ext : out    vl_logic;
        rxdata1_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak1_ext    : in     vl_logic;
        rxelecidle1_ext : in     vl_logic;
        rxpolarity1_ext : out    vl_logic;
        rxstatus1_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid1_ext    : in     vl_logic;
        txcompl1_ext    : out    vl_logic;
        txdata1_ext     : out    vl_logic_vector(7 downto 0);
        txdatak1_ext    : out    vl_logic;
        txelecidle1_ext : out    vl_logic;
        rxdata2_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak2_ext    : in     vl_logic;
        rxelecidle2_ext : in     vl_logic;
        rxpolarity2_ext : out    vl_logic;
        rxstatus2_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid2_ext    : in     vl_logic;
        txcompl2_ext    : out    vl_logic;
        txdata2_ext     : out    vl_logic_vector(7 downto 0);
        txdatak2_ext    : out    vl_logic;
        txelecidle2_ext : out    vl_logic;
        rxdata3_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak3_ext    : in     vl_logic;
        rxelecidle3_ext : in     vl_logic;
        rxpolarity3_ext : out    vl_logic;
        rxstatus3_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid3_ext    : in     vl_logic;
        txcompl3_ext    : out    vl_logic;
        txdata3_ext     : out    vl_logic_vector(7 downto 0);
        txdatak3_ext    : out    vl_logic;
        txelecidle3_ext : out    vl_logic;
        rxdata4_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak4_ext    : in     vl_logic;
        rxelecidle4_ext : in     vl_logic;
        rxpolarity4_ext : out    vl_logic;
        rxstatus4_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid4_ext    : in     vl_logic;
        txcompl4_ext    : out    vl_logic;
        txdata4_ext     : out    vl_logic_vector(7 downto 0);
        txdatak4_ext    : out    vl_logic;
        txelecidle4_ext : out    vl_logic;
        rxdata5_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak5_ext    : in     vl_logic;
        rxelecidle5_ext : in     vl_logic;
        rxpolarity5_ext : out    vl_logic;
        rxstatus5_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid5_ext    : in     vl_logic;
        txcompl5_ext    : out    vl_logic;
        txdata5_ext     : out    vl_logic_vector(7 downto 0);
        txdatak5_ext    : out    vl_logic;
        txelecidle5_ext : out    vl_logic;
        rxdata6_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak6_ext    : in     vl_logic;
        rxelecidle6_ext : in     vl_logic;
        rxpolarity6_ext : out    vl_logic;
        rxstatus6_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid6_ext    : in     vl_logic;
        txcompl6_ext    : out    vl_logic;
        txdata6_ext     : out    vl_logic_vector(7 downto 0);
        txdatak6_ext    : out    vl_logic;
        txelecidle6_ext : out    vl_logic;
        rxdata7_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak7_ext    : in     vl_logic;
        rxelecidle7_ext : in     vl_logic;
        rxpolarity7_ext : out    vl_logic;
        rxstatus7_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid7_ext    : in     vl_logic;
        txcompl7_ext    : out    vl_logic;
        txdata7_ext     : out    vl_logic_vector(7 downto 0);
        txdatak7_ext    : out    vl_logic;
        txelecidle7_ext : out    vl_logic;
        txdetectrx_ext  : out    vl_logic;
        cfg_devcsr      : out    vl_logic_vector(31 downto 0)
    );
end pcie_top;
