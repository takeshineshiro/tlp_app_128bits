library verilog;
use verilog.vl_types.all;
entity altpcietb_bfm_rpvar_64b_x8_pipen1b is
    port(
        app_int_sts     : in     vl_logic;
        app_msi_ack     : out    vl_logic;
        app_msi_req     : in     vl_logic;
        app_msi_tc      : in     vl_logic_vector(2 downto 0);
        cfg_busdev      : out    vl_logic_vector(12 downto 0);
        cfg_devcsr      : out    vl_logic_vector(31 downto 0);
        cfg_io_bas      : out    vl_logic_vector(19 downto 0);
        cfg_io_lim      : out    vl_logic_vector(19 downto 0);
        cfg_linkcsr     : out    vl_logic_vector(31 downto 0);
        cfg_msicsr      : out    vl_logic_vector(15 downto 0);
        cfg_np_bas      : out    vl_logic_vector(11 downto 0);
        cfg_np_lim      : out    vl_logic_vector(11 downto 0);
        cfg_pmcsr       : out    vl_logic_vector(31 downto 0);
        cfg_pr_bas      : out    vl_logic_vector(43 downto 0);
        cfg_pr_lim      : out    vl_logic_vector(43 downto 0);
        cfg_prmcsr      : out    vl_logic_vector(31 downto 0);
        cfg_rootcsr     : out    vl_logic_vector(31 downto 0);
        cfg_secbus      : out    vl_logic_vector(7 downto 0);
        cfg_seccsr      : out    vl_logic_vector(31 downto 0);
        cfg_slotcsr     : out    vl_logic_vector(31 downto 0);
        cfg_subbus      : out    vl_logic_vector(7 downto 0);
        cfg_tcvcmap     : out    vl_logic_vector(23 downto 0);
        coreclk_out     : out    vl_logic;
        cpl_err         : in     vl_logic_vector(2 downto 0);
        cpl_pending     : in     vl_logic;
        crst            : in     vl_logic;
        dlup_exit       : out    vl_logic;
        ep_clk250_in    : in     vl_logic;
        hotrst_exit     : out    vl_logic;
        l2_exit         : out    vl_logic;
        npor            : in     vl_logic;
        pclk_in         : in     vl_logic;
        phystatus0_ext  : in     vl_logic;
        phystatus1_ext  : in     vl_logic;
        phystatus2_ext  : in     vl_logic;
        phystatus3_ext  : in     vl_logic;
        phystatus4_ext  : in     vl_logic;
        phystatus5_ext  : in     vl_logic;
        phystatus6_ext  : in     vl_logic;
        phystatus7_ext  : in     vl_logic;
        pipe_mode       : in     vl_logic;
        pm_auxpwr       : in     vl_logic;
        pme_to_cr       : in     vl_logic;
        pme_to_sr       : out    vl_logic;
        powerdown0_ext  : out    vl_logic_vector(1 downto 0);
        powerdown1_ext  : out    vl_logic_vector(1 downto 0);
        powerdown2_ext  : out    vl_logic_vector(1 downto 0);
        powerdown3_ext  : out    vl_logic_vector(1 downto 0);
        powerdown4_ext  : out    vl_logic_vector(1 downto 0);
        powerdown5_ext  : out    vl_logic_vector(1 downto 0);
        powerdown6_ext  : out    vl_logic_vector(1 downto 0);
        powerdown7_ext  : out    vl_logic_vector(1 downto 0);
        rate_ext        : out    vl_logic;
        rx_abort0       : in     vl_logic;
        rx_abort1       : in     vl_logic;
        rx_abort2       : in     vl_logic;
        rx_abort3       : in     vl_logic;
        rx_ack0         : in     vl_logic;
        rx_ack1         : in     vl_logic;
        rx_ack2         : in     vl_logic;
        rx_ack3         : in     vl_logic;
        rx_be0          : out    vl_logic_vector(7 downto 0);
        rx_be1          : out    vl_logic_vector(7 downto 0);
        rx_be2          : out    vl_logic_vector(7 downto 0);
        rx_be3          : out    vl_logic_vector(7 downto 0);
        rx_data0        : out    vl_logic_vector(63 downto 0);
        rx_data1        : out    vl_logic_vector(63 downto 0);
        rx_data2        : out    vl_logic_vector(63 downto 0);
        rx_data3        : out    vl_logic_vector(63 downto 0);
        rx_desc0        : out    vl_logic_vector(135 downto 0);
        rx_desc1        : out    vl_logic_vector(135 downto 0);
        rx_desc2        : out    vl_logic_vector(135 downto 0);
        rx_desc3        : out    vl_logic_vector(135 downto 0);
        rx_dfr0         : out    vl_logic;
        rx_dfr1         : out    vl_logic;
        rx_dfr2         : out    vl_logic;
        rx_dfr3         : out    vl_logic;
        rx_dv0          : out    vl_logic;
        rx_dv1          : out    vl_logic;
        rx_dv2          : out    vl_logic;
        rx_dv3          : out    vl_logic;
        rx_in0          : in     vl_logic;
        rx_in1          : in     vl_logic;
        rx_in2          : in     vl_logic;
        rx_in3          : in     vl_logic;
        rx_in4          : in     vl_logic;
        rx_in5          : in     vl_logic;
        rx_in6          : in     vl_logic;
        rx_in7          : in     vl_logic;
        rx_mask0        : in     vl_logic;
        rx_mask1        : in     vl_logic;
        rx_mask2        : in     vl_logic;
        rx_mask3        : in     vl_logic;
        rx_req0         : out    vl_logic;
        rx_req1         : out    vl_logic;
        rx_req2         : out    vl_logic;
        rx_req3         : out    vl_logic;
        rx_retry0       : in     vl_logic;
        rx_retry1       : in     vl_logic;
        rx_retry2       : in     vl_logic;
        rx_retry3       : in     vl_logic;
        rx_ws0          : in     vl_logic;
        rx_ws1          : in     vl_logic;
        rx_ws2          : in     vl_logic;
        rx_ws3          : in     vl_logic;
        rxdata0_ext     : in     vl_logic_vector(7 downto 0);
        rxdata1_ext     : in     vl_logic_vector(7 downto 0);
        rxdata2_ext     : in     vl_logic_vector(7 downto 0);
        rxdata3_ext     : in     vl_logic_vector(7 downto 0);
        rxdata4_ext     : in     vl_logic_vector(7 downto 0);
        rxdata5_ext     : in     vl_logic_vector(7 downto 0);
        rxdata6_ext     : in     vl_logic_vector(7 downto 0);
        rxdata7_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak0_ext    : in     vl_logic;
        rxdatak1_ext    : in     vl_logic;
        rxdatak2_ext    : in     vl_logic;
        rxdatak3_ext    : in     vl_logic;
        rxdatak4_ext    : in     vl_logic;
        rxdatak5_ext    : in     vl_logic;
        rxdatak6_ext    : in     vl_logic;
        rxdatak7_ext    : in     vl_logic;
        rxelecidle0_ext : in     vl_logic;
        rxelecidle1_ext : in     vl_logic;
        rxelecidle2_ext : in     vl_logic;
        rxelecidle3_ext : in     vl_logic;
        rxelecidle4_ext : in     vl_logic;
        rxelecidle5_ext : in     vl_logic;
        rxelecidle6_ext : in     vl_logic;
        rxelecidle7_ext : in     vl_logic;
        rxpolarity0_ext : out    vl_logic;
        rxpolarity1_ext : out    vl_logic;
        rxpolarity2_ext : out    vl_logic;
        rxpolarity3_ext : out    vl_logic;
        rxpolarity4_ext : out    vl_logic;
        rxpolarity5_ext : out    vl_logic;
        rxpolarity6_ext : out    vl_logic;
        rxpolarity7_ext : out    vl_logic;
        rxstatus0_ext   : in     vl_logic_vector(2 downto 0);
        rxstatus1_ext   : in     vl_logic_vector(2 downto 0);
        rxstatus2_ext   : in     vl_logic_vector(2 downto 0);
        rxstatus3_ext   : in     vl_logic_vector(2 downto 0);
        rxstatus4_ext   : in     vl_logic_vector(2 downto 0);
        rxstatus5_ext   : in     vl_logic_vector(2 downto 0);
        rxstatus6_ext   : in     vl_logic_vector(2 downto 0);
        rxstatus7_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid0_ext    : in     vl_logic;
        rxvalid1_ext    : in     vl_logic;
        rxvalid2_ext    : in     vl_logic;
        rxvalid3_ext    : in     vl_logic;
        rxvalid4_ext    : in     vl_logic;
        rxvalid5_ext    : in     vl_logic;
        rxvalid6_ext    : in     vl_logic;
        rxvalid7_ext    : in     vl_logic;
        serr_out        : out    vl_logic;
        slotcap_in      : in     vl_logic_vector(6 downto 0);
        slotnum_in      : in     vl_logic_vector(12 downto 0);
        srst            : in     vl_logic;
        swdn_out        : out    vl_logic_vector(5 downto 0);
        test_in         : in     vl_logic_vector(31 downto 0);
        test_out        : out    vl_logic_vector(511 downto 0);
        tx_ack0         : out    vl_logic;
        tx_ack1         : out    vl_logic;
        tx_ack2         : out    vl_logic;
        tx_ack3         : out    vl_logic;
        tx_cred0        : out    vl_logic_vector(21 downto 0);
        tx_cred1        : out    vl_logic_vector(21 downto 0);
        tx_cred2        : out    vl_logic_vector(21 downto 0);
        tx_cred3        : out    vl_logic_vector(21 downto 0);
        tx_data0        : in     vl_logic_vector(63 downto 0);
        tx_data1        : in     vl_logic_vector(63 downto 0);
        tx_data2        : in     vl_logic_vector(63 downto 0);
        tx_data3        : in     vl_logic_vector(63 downto 0);
        tx_desc0        : in     vl_logic_vector(127 downto 0);
        tx_desc1        : in     vl_logic_vector(127 downto 0);
        tx_desc2        : in     vl_logic_vector(127 downto 0);
        tx_desc3        : in     vl_logic_vector(127 downto 0);
        tx_dfr0         : in     vl_logic;
        tx_dfr1         : in     vl_logic;
        tx_dfr2         : in     vl_logic;
        tx_dfr3         : in     vl_logic;
        tx_dv0          : in     vl_logic;
        tx_dv1          : in     vl_logic;
        tx_dv2          : in     vl_logic;
        tx_dv3          : in     vl_logic;
        tx_err0         : in     vl_logic;
        tx_err1         : in     vl_logic;
        tx_err2         : in     vl_logic;
        tx_err3         : in     vl_logic;
        tx_out0         : out    vl_logic;
        tx_out1         : out    vl_logic;
        tx_out2         : out    vl_logic;
        tx_out3         : out    vl_logic;
        tx_out4         : out    vl_logic;
        tx_out5         : out    vl_logic;
        tx_out6         : out    vl_logic;
        tx_out7         : out    vl_logic;
        tx_req0         : in     vl_logic;
        tx_req1         : in     vl_logic;
        tx_req2         : in     vl_logic;
        tx_req3         : in     vl_logic;
        tx_ws0          : out    vl_logic;
        tx_ws1          : out    vl_logic;
        tx_ws2          : out    vl_logic;
        tx_ws3          : out    vl_logic;
        txcompl0_ext    : out    vl_logic;
        txcompl1_ext    : out    vl_logic;
        txcompl2_ext    : out    vl_logic;
        txcompl3_ext    : out    vl_logic;
        txcompl4_ext    : out    vl_logic;
        txcompl5_ext    : out    vl_logic;
        txcompl6_ext    : out    vl_logic;
        txcompl7_ext    : out    vl_logic;
        txdata0_ext     : out    vl_logic_vector(7 downto 0);
        txdata1_ext     : out    vl_logic_vector(7 downto 0);
        txdata2_ext     : out    vl_logic_vector(7 downto 0);
        txdata3_ext     : out    vl_logic_vector(7 downto 0);
        txdata4_ext     : out    vl_logic_vector(7 downto 0);
        txdata5_ext     : out    vl_logic_vector(7 downto 0);
        txdata6_ext     : out    vl_logic_vector(7 downto 0);
        txdata7_ext     : out    vl_logic_vector(7 downto 0);
        txdatak0_ext    : out    vl_logic;
        txdatak1_ext    : out    vl_logic;
        txdatak2_ext    : out    vl_logic;
        txdatak3_ext    : out    vl_logic;
        txdatak4_ext    : out    vl_logic;
        txdatak5_ext    : out    vl_logic;
        txdatak6_ext    : out    vl_logic;
        txdatak7_ext    : out    vl_logic;
        txdetectrx0_ext : out    vl_logic;
        txdetectrx1_ext : out    vl_logic;
        txdetectrx2_ext : out    vl_logic;
        txdetectrx3_ext : out    vl_logic;
        txdetectrx4_ext : out    vl_logic;
        txdetectrx5_ext : out    vl_logic;
        txdetectrx6_ext : out    vl_logic;
        txdetectrx7_ext : out    vl_logic;
        txelecidle0_ext : out    vl_logic;
        txelecidle1_ext : out    vl_logic;
        txelecidle2_ext : out    vl_logic;
        txelecidle3_ext : out    vl_logic;
        txelecidle4_ext : out    vl_logic;
        txelecidle5_ext : out    vl_logic;
        txelecidle6_ext : out    vl_logic;
        txelecidle7_ext : out    vl_logic
    );
end altpcietb_bfm_rpvar_64b_x8_pipen1b;
