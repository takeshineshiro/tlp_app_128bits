library verilog;
use verilog.vl_types.all;
entity pcie_core is
    generic(
        PCIE_VENDOR_ID  : integer := 4466;
        PCIE_DEVICE_ID  : integer := 4;
        PCIE_VEVISION_ID: integer := 1
    );
    port(
        AvlClk_i        : in     vl_logic;
        CraAddress_i    : in     vl_logic_vector(11 downto 0);
        CraByteEnable_i : in     vl_logic_vector(3 downto 0);
        CraChipSelect_i : in     vl_logic;
        CraRead         : in     vl_logic;
        CraWrite        : in     vl_logic;
        CraWriteData_i  : in     vl_logic_vector(31 downto 0);
        Rstn_i          : in     vl_logic;
        RxmIrqNum_i     : in     vl_logic_vector(5 downto 0);
        RxmIrq_i        : in     vl_logic;
        RxmReadDataValid_i: in     vl_logic;
        RxmReadData_i   : in     vl_logic_vector(63 downto 0);
        RxmWaitRequest_i: in     vl_logic;
        TxsAddress_i    : in     vl_logic_vector(16 downto 0);
        TxsBurstCount_i : in     vl_logic_vector(9 downto 0);
        TxsByteEnable_i : in     vl_logic_vector(7 downto 0);
        TxsChipSelect_i : in     vl_logic;
        TxsRead_i       : in     vl_logic;
        TxsWriteData_i  : in     vl_logic_vector(63 downto 0);
        TxsWrite_i      : in     vl_logic;
        aer_msi_num     : in     vl_logic_vector(4 downto 0);
        app_int_sts     : in     vl_logic;
        app_msi_num     : in     vl_logic_vector(4 downto 0);
        app_msi_req     : in     vl_logic;
        app_msi_tc      : in     vl_logic_vector(2 downto 0);
        core_clk_in     : in     vl_logic;
        cpl_err         : in     vl_logic_vector(6 downto 0);
        cpl_pending     : in     vl_logic;
        crst            : in     vl_logic;
        hpg_ctrler      : in     vl_logic_vector(4 downto 0);
        lmi_addr        : in     vl_logic_vector(11 downto 0);
        lmi_din         : in     vl_logic_vector(31 downto 0);
        lmi_rden        : in     vl_logic;
        lmi_wren        : in     vl_logic;
        npor            : in     vl_logic;
        pclk_central    : in     vl_logic;
        pclk_ch0        : in     vl_logic;
        pex_msi_num     : in     vl_logic_vector(4 downto 0);
        pld_clk         : in     vl_logic;
        pll_fixed_clk   : in     vl_logic;
        pm_auxpwr       : in     vl_logic;
        pm_data         : in     vl_logic_vector(9 downto 0);
        pm_event        : in     vl_logic;
        pme_to_cr       : in     vl_logic;
        rc_areset       : in     vl_logic;
        rc_inclk_eq_125mhz: in     vl_logic;
        rc_pll_locked   : in     vl_logic;
        rc_rx_pll_locked_one: in     vl_logic;
        rx_st_mask0     : in     vl_logic;
        rx_st_ready0    : in     vl_logic;
        srst            : in     vl_logic;
        test_in         : in     vl_logic_vector(39 downto 0);
        tx_st_data0     : in     vl_logic_vector(63 downto 0);
        tx_st_data0_p1  : in     vl_logic_vector(63 downto 0);
        tx_st_eop0      : in     vl_logic;
        tx_st_eop0_p1   : in     vl_logic;
        tx_st_err0      : in     vl_logic;
        tx_st_sop0      : in     vl_logic;
        tx_st_sop0_p1   : in     vl_logic;
        tx_st_valid0    : in     vl_logic;
        phystatus0_ext  : in     vl_logic;
        rxdata0_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak0_ext    : in     vl_logic;
        rxelecidle0_ext : in     vl_logic;
        rxstatus0_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid0_ext    : in     vl_logic;
        phystatus1_ext  : in     vl_logic;
        rxdata1_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak1_ext    : in     vl_logic;
        rxelecidle1_ext : in     vl_logic;
        rxstatus1_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid1_ext    : in     vl_logic;
        phystatus2_ext  : in     vl_logic;
        rxdata2_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak2_ext    : in     vl_logic;
        rxelecidle2_ext : in     vl_logic;
        rxstatus2_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid2_ext    : in     vl_logic;
        phystatus3_ext  : in     vl_logic;
        rxdata3_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak3_ext    : in     vl_logic;
        rxelecidle3_ext : in     vl_logic;
        rxstatus3_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid3_ext    : in     vl_logic;
        phystatus4_ext  : in     vl_logic;
        rxdata4_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak4_ext    : in     vl_logic;
        rxelecidle4_ext : in     vl_logic;
        rxstatus4_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid4_ext    : in     vl_logic;
        phystatus5_ext  : in     vl_logic;
        rxdata5_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak5_ext    : in     vl_logic;
        rxelecidle5_ext : in     vl_logic;
        rxstatus5_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid5_ext    : in     vl_logic;
        phystatus6_ext  : in     vl_logic;
        rxdata6_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak6_ext    : in     vl_logic;
        rxelecidle6_ext : in     vl_logic;
        rxstatus6_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid6_ext    : in     vl_logic;
        phystatus7_ext  : in     vl_logic;
        rxdata7_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak7_ext    : in     vl_logic;
        rxelecidle7_ext : in     vl_logic;
        rxstatus7_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid7_ext    : in     vl_logic;
        CraIrq_o        : out    vl_logic;
        CraReadData_o   : out    vl_logic_vector(31 downto 0);
        CraWaitRequest_o: out    vl_logic;
        RxmAddress_o    : out    vl_logic_vector(31 downto 0);
        RxmBurstCount_o : out    vl_logic_vector(9 downto 0);
        RxmByteEnable_o : out    vl_logic_vector(7 downto 0);
        RxmRead_o       : out    vl_logic;
        RxmWriteData_o  : out    vl_logic_vector(63 downto 0);
        RxmWrite_o      : out    vl_logic;
        TxsReadDataValid_o: out    vl_logic;
        TxsReadData_o   : out    vl_logic_vector(63 downto 0);
        TxsWaitRequest_o: out    vl_logic;
        app_int_ack     : out    vl_logic;
        app_msi_ack     : out    vl_logic;
        avs_pcie_reconfig_readdata: out    vl_logic_vector(15 downto 0);
        avs_pcie_reconfig_readdatavalid: out    vl_logic;
        avs_pcie_reconfig_waitrequest: out    vl_logic;
        core_clk_out    : out    vl_logic;
        derr_cor_ext_rcv0: out    vl_logic;
        derr_cor_ext_rpl: out    vl_logic;
        derr_rpl        : out    vl_logic;
        dl_ltssm        : out    vl_logic_vector(4 downto 0);
        dlup_exit       : out    vl_logic;
        eidle_infer_sel : out    vl_logic_vector(23 downto 0);
        ev_128ns        : out    vl_logic;
        ev_1us          : out    vl_logic;
        hip_extraclkout : out    vl_logic_vector(1 downto 0);
        hotrst_exit     : out    vl_logic;
        int_status      : out    vl_logic_vector(3 downto 0);
        l2_exit         : out    vl_logic;
        lane_act        : out    vl_logic_vector(3 downto 0);
        lmi_ack         : out    vl_logic;
        lmi_dout        : out    vl_logic_vector(31 downto 0);
        npd_alloc_1cred_vc0: out    vl_logic;
        npd_cred_vio_vc0: out    vl_logic;
        nph_alloc_1cred_vc0: out    vl_logic;
        nph_cred_vio_vc0: out    vl_logic;
        pme_to_sr       : out    vl_logic;
        r2c_err0        : out    vl_logic;
        rate_ext        : out    vl_logic;
        rc_gxb_powerdown: out    vl_logic;
        rc_rx_analogreset: out    vl_logic;
        rc_rx_digitalreset: out    vl_logic;
        rc_tx_digitalreset: out    vl_logic;
        reset_status    : out    vl_logic;
        rx_fifo_empty0  : out    vl_logic;
        rx_fifo_full0   : out    vl_logic;
        rx_st_bardec0   : out    vl_logic_vector(7 downto 0);
        rx_st_be0       : out    vl_logic_vector(7 downto 0);
        rx_st_be0_p1    : out    vl_logic_vector(7 downto 0);
        rx_st_data0     : out    vl_logic_vector(63 downto 0);
        rx_st_data0_p1  : out    vl_logic_vector(63 downto 0);
        rx_st_eop0      : out    vl_logic;
        rx_st_eop0_p1   : out    vl_logic;
        rx_st_err0      : out    vl_logic;
        rx_st_sop0      : out    vl_logic;
        rx_st_sop0_p1   : out    vl_logic;
        rx_st_valid0    : out    vl_logic;
        serr_out        : out    vl_logic;
        suc_spd_neg     : out    vl_logic;
        swdn_wake       : out    vl_logic;
        swup_hotrst     : out    vl_logic;
        test_out        : out    vl_logic_vector(63 downto 0);
        tl_cfg_add      : out    vl_logic_vector(3 downto 0);
        tl_cfg_ctl      : out    vl_logic_vector(31 downto 0);
        tl_cfg_ctl_wr   : out    vl_logic;
        tl_cfg_sts      : out    vl_logic_vector(52 downto 0);
        tl_cfg_sts_wr   : out    vl_logic;
        tx_cred0        : out    vl_logic_vector(35 downto 0);
        tx_deemph       : out    vl_logic_vector(7 downto 0);
        tx_fifo_empty0  : out    vl_logic;
        tx_fifo_full0   : out    vl_logic;
        tx_fifo_rdptr0  : out    vl_logic_vector(3 downto 0);
        tx_fifo_wrptr0  : out    vl_logic_vector(3 downto 0);
        tx_margin       : out    vl_logic_vector(23 downto 0);
        tx_st_ready0    : out    vl_logic;
        use_pcie_reconfig: out    vl_logic;
        wake_oen        : out    vl_logic;
        powerdown0_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity0_ext : out    vl_logic;
        txcompl0_ext    : out    vl_logic;
        txdata0_ext     : out    vl_logic_vector(7 downto 0);
        txdatak0_ext    : out    vl_logic;
        txdetectrx0_ext : out    vl_logic;
        txelecidle0_ext : out    vl_logic;
        powerdown1_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity1_ext : out    vl_logic;
        txcompl1_ext    : out    vl_logic;
        txdata1_ext     : out    vl_logic_vector(7 downto 0);
        txdatak1_ext    : out    vl_logic;
        txdetectrx1_ext : out    vl_logic;
        txelecidle1_ext : out    vl_logic;
        powerdown2_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity2_ext : out    vl_logic;
        txcompl2_ext    : out    vl_logic;
        txdata2_ext     : out    vl_logic_vector(7 downto 0);
        txdatak2_ext    : out    vl_logic;
        txdetectrx2_ext : out    vl_logic;
        txelecidle2_ext : out    vl_logic;
        powerdown3_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity3_ext : out    vl_logic;
        txcompl3_ext    : out    vl_logic;
        txdata3_ext     : out    vl_logic_vector(7 downto 0);
        txdatak3_ext    : out    vl_logic;
        txdetectrx3_ext : out    vl_logic;
        txelecidle3_ext : out    vl_logic;
        powerdown4_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity4_ext : out    vl_logic;
        txcompl4_ext    : out    vl_logic;
        txdata4_ext     : out    vl_logic_vector(7 downto 0);
        txdatak4_ext    : out    vl_logic;
        txdetectrx4_ext : out    vl_logic;
        txelecidle4_ext : out    vl_logic;
        powerdown5_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity5_ext : out    vl_logic;
        txcompl5_ext    : out    vl_logic;
        txdata5_ext     : out    vl_logic_vector(7 downto 0);
        txdatak5_ext    : out    vl_logic;
        txdetectrx5_ext : out    vl_logic;
        txelecidle5_ext : out    vl_logic;
        powerdown6_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity6_ext : out    vl_logic;
        txcompl6_ext    : out    vl_logic;
        txdata6_ext     : out    vl_logic_vector(7 downto 0);
        txdatak6_ext    : out    vl_logic;
        txdetectrx6_ext : out    vl_logic;
        txelecidle6_ext : out    vl_logic;
        powerdown7_ext  : out    vl_logic_vector(1 downto 0);
        rxpolarity7_ext : out    vl_logic;
        txcompl7_ext    : out    vl_logic;
        txdata7_ext     : out    vl_logic_vector(7 downto 0);
        txdatak7_ext    : out    vl_logic;
        txdetectrx7_ext : out    vl_logic;
        txelecidle7_ext : out    vl_logic
    );
end pcie_core;
