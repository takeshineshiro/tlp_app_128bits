library verilog;
use verilog.vl_types.all;
entity altpcietb_bfm_vc_intf is
    generic(
        VC_NUM          : integer := 0;
        DISABLE_RX_BE_CHECK: integer := 1;
        RP_PRI_BUS_NUM  : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RP_PRI_DEV_NUM  : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        SHMEM_ADDR_WIDTH: integer := 21;
        EBFM_BAR_M64_MIN: vl_logic_vector(63 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EBFM_NUM_VC     : integer := 4;
        EBFM_NUM_TAG    : integer := 32;
        EBFM_MSG_DEBUG  : integer := 0;
        EBFM_MSG_INFO   : integer := 1;
        EBFM_MSG_WARNING: integer := 2;
        EBFM_MSG_ERROR_INFO: integer := 3;
        EBFM_MSG_ERROR_CONTINUE: integer := 4;
        EBFM_MSG_ERROR_FATAL: integer := 101;
        EBFM_MSG_ERROR_FATAL_TB_ERR: integer := 102;
        EBFM_MSG_MAX_LEN: integer := 100;
        SHMEM_FILL_ZERO : integer := 0;
        SHMEM_FILL_BYTE_INC: integer := 1;
        SHMEM_FILL_WORD_INC: integer := 2;
        SHMEM_FILL_DWORD_INC: integer := 4;
        SHMEM_FILL_QWORD_INC: integer := 8;
        SHMEM_FILL_ONE  : integer := 15;
        BAR_TABLE_SIZE  : integer := 64;
        SCR_SIZE        : integer := 64;
        NUM_PS_TO_WAIT  : integer := 8000;
        RXST_IDLE       : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        RXST_DESC_ACK   : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        RXST_DATA_WRITE : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        RXST_DATA_NONP_WRITE: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        RXST_DATA_COMPL : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        RXST_NONP_REQ   : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1);
        TXST_IDLE       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        TXST_DESC       : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        TXST_DATA       : vl_logic_vector(1 downto 0) := (Hi1, Hi0)
    );
    port(
        clk_in          : in     vl_logic;
        rstn            : in     vl_logic;
        rx_req          : in     vl_logic;
        rx_ack          : out    vl_logic;
        rx_abort        : out    vl_logic;
        rx_retry        : out    vl_logic;
        rx_mask         : out    vl_logic;
        rx_desc         : in     vl_logic_vector(135 downto 0);
        rx_ws           : out    vl_logic;
        rx_data         : in     vl_logic_vector(63 downto 0);
        rx_be           : in     vl_logic_vector(7 downto 0);
        rx_dv           : in     vl_logic;
        rx_dfr          : in     vl_logic;
        tx_cred         : in     vl_logic_vector(21 downto 0);
        tx_req          : out    vl_logic;
        tx_desc         : out    vl_logic_vector(127 downto 0);
        tx_ack          : in     vl_logic;
        tx_dfr          : out    vl_logic;
        tx_data         : out    vl_logic_vector(63 downto 0);
        tx_dv           : out    vl_logic;
        tx_err          : out    vl_logic;
        tx_ws           : in     vl_logic;
        cfg_io_bas      : in     vl_logic_vector(19 downto 0);
        cfg_np_bas      : in     vl_logic_vector(11 downto 0);
        cfg_pr_bas      : in     vl_logic_vector(43 downto 0)
    );
    attribute RP_PRI_BUS_NUM_mti_vect_attrib : integer;
    attribute RP_PRI_BUS_NUM_mti_vect_attrib of RP_PRI_BUS_NUM : constant is 0;
    attribute RP_PRI_DEV_NUM_mti_vect_attrib : integer;
    attribute RP_PRI_DEV_NUM_mti_vect_attrib of RP_PRI_DEV_NUM : constant is 0;
    attribute EBFM_BAR_M64_MIN_mti_vect_attrib : integer;
    attribute EBFM_BAR_M64_MIN_mti_vect_attrib of EBFM_BAR_M64_MIN : constant is 0;
    attribute RXST_IDLE_mti_vect_attrib : integer;
    attribute RXST_IDLE_mti_vect_attrib of RXST_IDLE : constant is 0;
    attribute RXST_DESC_ACK_mti_vect_attrib : integer;
    attribute RXST_DESC_ACK_mti_vect_attrib of RXST_DESC_ACK : constant is 1;
    attribute RXST_DATA_WRITE_mti_vect_attrib : integer;
    attribute RXST_DATA_WRITE_mti_vect_attrib of RXST_DATA_WRITE : constant is 2;
    attribute RXST_DATA_NONP_WRITE_mti_vect_attrib : integer;
    attribute RXST_DATA_NONP_WRITE_mti_vect_attrib of RXST_DATA_NONP_WRITE : constant is 3;
    attribute RXST_DATA_COMPL_mti_vect_attrib : integer;
    attribute RXST_DATA_COMPL_mti_vect_attrib of RXST_DATA_COMPL : constant is 4;
    attribute RXST_NONP_REQ_mti_vect_attrib : integer;
    attribute RXST_NONP_REQ_mti_vect_attrib of RXST_NONP_REQ : constant is 5;
    attribute TXST_IDLE_mti_vect_attrib : integer;
    attribute TXST_IDLE_mti_vect_attrib of TXST_IDLE : constant is 0;
    attribute TXST_DESC_mti_vect_attrib : integer;
    attribute TXST_DESC_mti_vect_attrib of TXST_DESC : constant is 1;
    attribute TXST_DATA_mti_vect_attrib : integer;
    attribute TXST_DATA_mti_vect_attrib of TXST_DATA : constant is 2;
end altpcietb_bfm_vc_intf;
