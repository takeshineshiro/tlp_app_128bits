library verilog;
use verilog.vl_types.all;
entity ict106_si_transactor is
    generic(
        C_MAX_M         : integer := 16;
        C_NUM_ADDR_RANGES: integer := 16;
        C_FAMILY        : string  := "none";
        C_SI            : integer := 0;
        C_DIR           : integer := 0;
        C_NUM_M         : integer := 2;
        C_NUM_M_LOG     : integer := 1;
        C_ACCEPTANCE    : integer := 1;
        C_ACCEPTANCE_LOG: integer := 0;
        C_ID_WIDTH      : integer := 1;
        C_ADDR_WIDTH    : integer := 32;
        C_AMESG_WIDTH   : integer := 1;
        C_RMESG_WIDTH   : integer := 1;
        C_THREAD_ID_WIDTH: integer := 0;
        C_BASE_ID       : vl_logic_vector(63 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        C_HIGH_ID       : vl_logic_vector(63 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        C_IS_INTERCONNECT: integer := 0;
        C_TARGET_QUAL   : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        C_SINGLE_THREAD : integer := 0;
        C_RANGE_CHECK   : integer := 0;
        C_ADDR_DECODE   : integer := 0;
        C_DEBUG         : integer := 1;
        C_MAX_DEBUG_THREADS: integer := 1
    );
    port(
        ACLK            : in     vl_logic;
        ARESET          : in     vl_logic;
        S_AID           : in     vl_logic_vector;
        S_AADDR         : in     vl_logic_vector;
        S_ALEN          : in     vl_logic_vector(7 downto 0);
        S_ASIZE         : in     vl_logic_vector(2 downto 0);
        S_ABURST        : in     vl_logic_vector(1 downto 0);
        S_ALOCK         : in     vl_logic_vector(1 downto 0);
        S_APROT         : in     vl_logic_vector(2 downto 0);
        S_AMESG         : in     vl_logic_vector;
        S_AVALID        : in     vl_logic;
        S_AREADY        : out    vl_logic;
        M_AID           : out    vl_logic_vector;
        M_AADDR         : out    vl_logic_vector;
        M_ALEN          : out    vl_logic_vector(7 downto 0);
        M_ASIZE         : out    vl_logic_vector(2 downto 0);
        M_ALOCK         : out    vl_logic_vector(1 downto 0);
        M_APROT         : out    vl_logic_vector(2 downto 0);
        M_AREGION       : out    vl_logic_vector(3 downto 0);
        M_AMESG         : out    vl_logic_vector;
        M_ATARGET_HOT   : out    vl_logic_vector;
        M_ATARGET_ENC   : out    vl_logic_vector;
        M_AERROR        : out    vl_logic_vector(7 downto 0);
        M_AVALID_QUAL   : out    vl_logic;
        M_AVALID        : out    vl_logic;
        M_AREADY        : in     vl_logic;
        S_RID           : out    vl_logic_vector;
        S_RMESG         : out    vl_logic_vector;
        S_RLAST         : out    vl_logic;
        S_RVALID        : out    vl_logic;
        S_RREADY        : in     vl_logic;
        M_RID           : in     vl_logic_vector;
        M_RMESG         : in     vl_logic_vector;
        M_RLAST         : in     vl_logic_vector;
        M_RVALID        : in     vl_logic_vector;
        M_RREADY        : out    vl_logic_vector;
        M_RTARGET       : in     vl_logic_vector;
        DEBUG_A_TRANS_SEQ: in     vl_logic_vector(7 downto 0);
        DEBUG_ACCEPT_CNT: out    vl_logic_vector;
        DEBUG_ACTIVE_THREAD: out    vl_logic_vector(15 downto 0);
        DEBUG_ACTIVE_TARGET: out    vl_logic_vector;
        DEBUG_ACTIVE_REGION: out    vl_logic_vector;
        DEBUG_R_BEAT_CNT: out    vl_logic_vector;
        DEBUG_R_TRANS_SEQ: out    vl_logic_vector;
        DEBUG_TRANS_QUAL: out    vl_logic_vector
    );
    attribute C_BASE_ID_mti_vect_attrib : integer;
    attribute C_BASE_ID_mti_vect_attrib of C_BASE_ID : constant is -1;
    attribute C_HIGH_ID_mti_vect_attrib : integer;
    attribute C_HIGH_ID_mti_vect_attrib of C_HIGH_ID : constant is 0;
    attribute C_TARGET_QUAL_mti_vect_attrib : integer;
    attribute C_TARGET_QUAL_mti_vect_attrib of C_TARGET_QUAL : constant is -1;
end ict106_si_transactor;
