library verilog;
use verilog.vl_types.all;
entity top is
    generic(
        AXI_DATA_WIDTH  : integer := 64;
        AXI_ADDR_WIDTH  : integer := 32;
        USER_WIDTH_RX   : integer := 22;
        USER_WIDTH_TX   : integer := 4;
        AXI_ID_WIDTH    : integer := 4;
        C_PIPE_MODE     : integer := 0;
        C_NO_OF_LANES   : integer := 8
    );
    port(
        pcie_rstn       : in     vl_logic;
        refclk          : in     vl_logic;
        free_100MHz     : in     vl_logic;
        core_clk_out    : out    vl_logic;
        linkdown        : out    vl_logic;
        fan_con         : out    vl_logic;
        pci_exp_rxp     : in     vl_logic_vector;
        pci_exp_txp     : out    vl_logic_vector;
        test_in         : in     vl_logic_vector(39 downto 0);
        test_out_icm    : out    vl_logic_vector(8 downto 0);
        phystatus_ext   : in     vl_logic;
        powerdown_ext   : out    vl_logic_vector(1 downto 0);
        rate_ext        : out    vl_logic;
        pclk_in         : in     vl_logic;
        clk250_out      : out    vl_logic;
        clk500_out      : out    vl_logic;
        rxdata0_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak0_ext    : in     vl_logic;
        rxelecidle0_ext : in     vl_logic;
        rxpolarity0_ext : out    vl_logic;
        rxstatus0_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid0_ext    : in     vl_logic;
        txcompl0_ext    : out    vl_logic;
        txdata0_ext     : out    vl_logic_vector(7 downto 0);
        txdatak0_ext    : out    vl_logic;
        txelecidle0_ext : out    vl_logic;
        rxdata1_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak1_ext    : in     vl_logic;
        rxelecidle1_ext : in     vl_logic;
        rxpolarity1_ext : out    vl_logic;
        rxstatus1_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid1_ext    : in     vl_logic;
        txcompl1_ext    : out    vl_logic;
        txdata1_ext     : out    vl_logic_vector(7 downto 0);
        txdatak1_ext    : out    vl_logic;
        txelecidle1_ext : out    vl_logic;
        rxdata2_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak2_ext    : in     vl_logic;
        rxelecidle2_ext : in     vl_logic;
        rxpolarity2_ext : out    vl_logic;
        rxstatus2_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid2_ext    : in     vl_logic;
        txcompl2_ext    : out    vl_logic;
        txdata2_ext     : out    vl_logic_vector(7 downto 0);
        txdatak2_ext    : out    vl_logic;
        txelecidle2_ext : out    vl_logic;
        rxdata3_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak3_ext    : in     vl_logic;
        rxelecidle3_ext : in     vl_logic;
        rxpolarity3_ext : out    vl_logic;
        rxstatus3_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid3_ext    : in     vl_logic;
        txcompl3_ext    : out    vl_logic;
        txdata3_ext     : out    vl_logic_vector(7 downto 0);
        txdatak3_ext    : out    vl_logic;
        txelecidle3_ext : out    vl_logic;
        rxdata4_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak4_ext    : in     vl_logic;
        rxelecidle4_ext : in     vl_logic;
        rxpolarity4_ext : out    vl_logic;
        rxstatus4_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid4_ext    : in     vl_logic;
        txcompl4_ext    : out    vl_logic;
        txdata4_ext     : out    vl_logic_vector(7 downto 0);
        txdatak4_ext    : out    vl_logic;
        txelecidle4_ext : out    vl_logic;
        rxdata5_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak5_ext    : in     vl_logic;
        rxelecidle5_ext : in     vl_logic;
        rxpolarity5_ext : out    vl_logic;
        rxstatus5_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid5_ext    : in     vl_logic;
        txcompl5_ext    : out    vl_logic;
        txdata5_ext     : out    vl_logic_vector(7 downto 0);
        txdatak5_ext    : out    vl_logic;
        txelecidle5_ext : out    vl_logic;
        rxdata6_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak6_ext    : in     vl_logic;
        rxelecidle6_ext : in     vl_logic;
        rxpolarity6_ext : out    vl_logic;
        rxstatus6_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid6_ext    : in     vl_logic;
        txcompl6_ext    : out    vl_logic;
        txdata6_ext     : out    vl_logic_vector(7 downto 0);
        txdatak6_ext    : out    vl_logic;
        txelecidle6_ext : out    vl_logic;
        rxdata7_ext     : in     vl_logic_vector(7 downto 0);
        rxdatak7_ext    : in     vl_logic;
        rxelecidle7_ext : in     vl_logic;
        rxpolarity7_ext : out    vl_logic;
        rxstatus7_ext   : in     vl_logic_vector(2 downto 0);
        rxvalid7_ext    : in     vl_logic;
        txcompl7_ext    : out    vl_logic;
        txdata7_ext     : out    vl_logic_vector(7 downto 0);
        txdatak7_ext    : out    vl_logic;
        txelecidle7_ext : out    vl_logic;
        txdetectrx_ext  : out    vl_logic
    );
end top;
